`timescale 1ns / 1ps
module Multiplier_32(
    input [31:0] A,
    input [31:0] B,
    output [63:0] product
);
wire [63:0] p0;
wire [63:0] p1;
wire [63:0] p2;
wire [63:0] p3;
wire [63:0] p4;
wire [63:0] p5;
wire [63:0] p6;
wire [63:0] p7;
wire [63:0] p8;
wire [63:0] p9;
wire [63:0] p10;
wire [63:0] p11;
wire [63:0] p12;
wire [63:0] p13;
wire [63:0] p14;
wire [63:0] p15;
wire c0,c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15;
booth b0(	
	.y2(B[1]),
	.y1(B[0]),
	.y0(0),
	.X({{32{A[31]}},A[31:0]}),
	.p(p0),
	.c(c0)
);
booth b1(
	.y2(B[3]),
	.y1(B[2]),
	.y0(B[1]),
	.X({{30{A[31]}},A[31:0],2'b0}),
	.p(p1),
	.c(c1)
);
booth b2(
	.y2(B[5]),
	.y1(B[4]),
	.y0(B[3]),
	.X({{28{A[31]}},A[31:0],4'b0}),
	.p(p2),
	.c(c2)
);
booth b3(
	.y2(B[7]),
	.y1(B[6]),
	.y0(B[5]),
	.X({{26{A[31]}},A[31:0],6'b0}),
	.p(p3),
	.c(c3)
);
booth b4(
	.y2(B[9]),
	.y1(B[8]),
	.y0(B[7]),
	.X({{24{A[31]}},A[31:0],8'b0}),
	.p(p4),
	.c(c4)
);
booth b5(
	.y2(B[11]),
	.y1(B[10]),
	.y0(B[9]),
	.X({{22{A[31]}},A[31:0],10'b0}),
	.p(p5),
	.c(c5)
);
booth b6(
	.y2(B[13]),
	.y1(B[12]),
	.y0(B[11]),
	.X({{20{A[31]}},A[31:0],12'b0}),
	.p(p6),
	.c(c6)
);
booth b7(
	.y2(B[15]),
	.y1(B[14]),
	.y0(B[13]),
	.X({{18{A[31]}},A[31:0],14'b0}),
	.p(p7),
	.c(c7)
);
booth b8(
	.y2(B[17]),
	.y1(B[16]),
	.y0(B[15]),
	.X({{16{A[31]}},A[31:0],16'b0}),
	.p(p8),
	.c(c8)
);
booth b9(
	.y2(B[19]),
	.y1(B[18]),
	.y0(B[17]),
	.X({{14{A[31]}},A[31:0],18'b0}),
	.p(p9),
	.c(c9)
);
booth b10(
	.y2(B[21]),
	.y1(B[20]),
	.y0(B[19]),
	.X({{12{A[31]}},A[31:0],20'b0}),
	.p(p10),
	.c(c10)
);
booth b11(
	.y2(B[23]),
	.y1(B[22]),
	.y0(B[21]),
	.X({{10{A[31]}},A[31:0],22'b0}),
	.p(p11),
	.c(c11)
);
booth b12(
	.y2(B[25]),
	.y1(B[24]),
	.y0(B[23]),
	.X({{8{A[31]}},A[31:0],24'b0}),
	.p(p12),
	.c(c12)
);
booth b13(
	.y2(B[27]),
	.y1(B[26]),
	.y0(B[25]),
	.X({{6{A[31]}},A[31:0],26'b0}),
	.p(p13),
	.c(c13)
);
booth b14(
	.y2(B[29]),
	.y1(B[28]),
	.y0(B[27]),
	.X({{4{A[31]}},A[31:0],28'b0}),
	.p(p14),
	.c(c14)
);
booth b15(
	.y2(B[31]),
	.y1(B[30]),
	.y0(B[29]),
	.X({{2{A[31]}},A[31:0],30'b0}),
	.p(p15),
	.c(c15)
);

wire cout0_0,cout0_1,cout0_2,cout0_3,cout0_4,cout0_5,cout0_6,cout0_7,cout0_8,cout0_9,cout0_10,cout0_11,cout0_12,cout0_13,cout1_0,cout1_1,cout1_2,cout1_3,cout1_4,cout1_5,cout1_6,cout1_7,cout1_8,cout1_9,cout1_10,cout1_11,cout1_12,cout1_13,cout2_0,cout2_1,cout2_2,cout2_3,cout2_4,cout2_5,cout2_6,cout2_7,cout2_8,cout2_9,cout2_10,cout2_11,cout2_12,cout2_13,cout3_0,cout3_1,cout3_2,cout3_3,cout3_4,cout3_5,cout3_6,cout3_7,cout3_8,cout3_9,cout3_10,cout3_11,cout3_12,cout3_13,cout4_0,cout4_1,cout4_2,cout4_3,cout4_4,cout4_5,cout4_6,cout4_7,cout4_8,cout4_9,cout4_10,cout4_11,cout4_12,cout4_13,cout5_0,cout5_1,cout5_2,cout5_3,cout5_4,cout5_5,cout5_6,cout5_7,cout5_8,cout5_9,cout5_10,cout5_11,cout5_12,cout5_13,cout6_0,cout6_1,cout6_2,cout6_3,cout6_4,cout6_5,cout6_6,cout6_7,cout6_8,cout6_9,cout6_10,cout6_11,cout6_12,cout6_13,cout7_0,cout7_1,cout7_2,cout7_3,cout7_4,cout7_5,cout7_6,cout7_7,cout7_8,cout7_9,cout7_10,cout7_11,cout7_12,cout7_13,cout8_0,cout8_1,cout8_2,cout8_3,cout8_4,cout8_5,cout8_6,cout8_7,cout8_8,cout8_9,cout8_10,cout8_11,cout8_12,cout8_13,cout9_0,cout9_1,cout9_2,cout9_3,cout9_4,cout9_5,cout9_6,cout9_7,cout9_8,cout9_9,cout9_10,cout9_11,cout9_12,cout9_13,cout10_0,cout10_1,cout10_2,cout10_3,cout10_4,cout10_5,cout10_6,cout10_7,cout10_8,cout10_9,cout10_10,cout10_11,cout10_12,cout10_13,cout11_0,cout11_1,cout11_2,cout11_3,cout11_4,cout11_5,cout11_6,cout11_7,cout11_8,cout11_9,cout11_10,cout11_11,cout11_12,cout11_13,cout12_0,cout12_1,cout12_2,cout12_3,cout12_4,cout12_5,cout12_6,cout12_7,cout12_8,cout12_9,cout12_10,cout12_11,cout12_12,cout12_13,cout13_0,cout13_1,cout13_2,cout13_3,cout13_4,cout13_5,cout13_6,cout13_7,cout13_8,cout13_9,cout13_10,cout13_11,cout13_12,cout13_13,cout14_0,cout14_1,cout14_2,cout14_3,cout14_4,cout14_5,cout14_6,cout14_7,cout14_8,cout14_9,cout14_10,cout14_11,cout14_12,cout14_13,cout15_0,cout15_1,cout15_2,cout15_3,cout15_4,cout15_5,cout15_6,cout15_7,cout15_8,cout15_9,cout15_10,cout15_11,cout15_12,cout15_13,cout16_0,cout16_1,cout16_2,cout16_3,cout16_4,cout16_5,cout16_6,cout16_7,cout16_8,cout16_9,cout16_10,cout16_11,cout16_12,cout16_13,cout17_0,cout17_1,cout17_2,cout17_3,cout17_4,cout17_5,cout17_6,cout17_7,cout17_8,cout17_9,cout17_10,cout17_11,cout17_12,cout17_13,cout18_0,cout18_1,cout18_2,cout18_3,cout18_4,cout18_5,cout18_6,cout18_7,cout18_8,cout18_9,cout18_10,cout18_11,cout18_12,cout18_13,cout19_0,cout19_1,cout19_2,cout19_3,cout19_4,cout19_5,cout19_6,cout19_7,cout19_8,cout19_9,cout19_10,cout19_11,cout19_12,cout19_13,cout20_0,cout20_1,cout20_2,cout20_3,cout20_4,cout20_5,cout20_6,cout20_7,cout20_8,cout20_9,cout20_10,cout20_11,cout20_12,cout20_13,cout21_0,cout21_1,cout21_2,cout21_3,cout21_4,cout21_5,cout21_6,cout21_7,cout21_8,cout21_9,cout21_10,cout21_11,cout21_12,cout21_13,cout22_0,cout22_1,cout22_2,cout22_3,cout22_4,cout22_5,cout22_6,cout22_7,cout22_8,cout22_9,cout22_10,cout22_11,cout22_12,cout22_13,cout23_0,cout23_1,cout23_2,cout23_3,cout23_4,cout23_5,cout23_6,cout23_7,cout23_8,cout23_9,cout23_10,cout23_11,cout23_12,cout23_13,cout24_0,cout24_1,cout24_2,cout24_3,cout24_4,cout24_5,cout24_6,cout24_7,cout24_8,cout24_9,cout24_10,cout24_11,cout24_12,cout24_13,cout25_0,cout25_1,cout25_2,cout25_3,cout25_4,cout25_5,cout25_6,cout25_7,cout25_8,cout25_9,cout25_10,cout25_11,cout25_12,cout25_13,cout26_0,cout26_1,cout26_2,cout26_3,cout26_4,cout26_5,cout26_6,cout26_7,cout26_8,cout26_9,cout26_10,cout26_11,cout26_12,cout26_13,cout27_0,cout27_1,cout27_2,cout27_3,cout27_4,cout27_5,cout27_6,cout27_7,cout27_8,cout27_9,cout27_10,cout27_11,cout27_12,cout27_13,cout28_0,cout28_1,cout28_2,cout28_3,cout28_4,cout28_5,cout28_6,cout28_7,cout28_8,cout28_9,cout28_10,cout28_11,cout28_12,cout28_13,cout29_0,cout29_1,cout29_2,cout29_3,cout29_4,cout29_5,cout29_6,cout29_7,cout29_8,cout29_9,cout29_10,cout29_11,cout29_12,cout29_13,cout30_0,cout30_1,cout30_2,cout30_3,cout30_4,cout30_5,cout30_6,cout30_7,cout30_8,cout30_9,cout30_10,cout30_11,cout30_12,cout30_13,cout31_0,cout31_1,cout31_2,cout31_3,cout31_4,cout31_5,cout31_6,cout31_7,cout31_8,cout31_9,cout31_10,cout31_11,cout31_12,cout31_13,cout32_0,cout32_1,cout32_2,cout32_3,cout32_4,cout32_5,cout32_6,cout32_7,cout32_8,cout32_9,cout32_10,cout32_11,cout32_12,cout32_13,cout33_0,cout33_1,cout33_2,cout33_3,cout33_4,cout33_5,cout33_6,cout33_7,cout33_8,cout33_9,cout33_10,cout33_11,cout33_12,cout33_13,cout34_0,cout34_1,cout34_2,cout34_3,cout34_4,cout34_5,cout34_6,cout34_7,cout34_8,cout34_9,cout34_10,cout34_11,cout34_12,cout34_13,cout35_0,cout35_1,cout35_2,cout35_3,cout35_4,cout35_5,cout35_6,cout35_7,cout35_8,cout35_9,cout35_10,cout35_11,cout35_12,cout35_13,cout36_0,cout36_1,cout36_2,cout36_3,cout36_4,cout36_5,cout36_6,cout36_7,cout36_8,cout36_9,cout36_10,cout36_11,cout36_12,cout36_13,cout37_0,cout37_1,cout37_2,cout37_3,cout37_4,cout37_5,cout37_6,cout37_7,cout37_8,cout37_9,cout37_10,cout37_11,cout37_12,cout37_13,cout38_0,cout38_1,cout38_2,cout38_3,cout38_4,cout38_5,cout38_6,cout38_7,cout38_8,cout38_9,cout38_10,cout38_11,cout38_12,cout38_13,cout39_0,cout39_1,cout39_2,cout39_3,cout39_4,cout39_5,cout39_6,cout39_7,cout39_8,cout39_9,cout39_10,cout39_11,cout39_12,cout39_13,cout40_0,cout40_1,cout40_2,cout40_3,cout40_4,cout40_5,cout40_6,cout40_7,cout40_8,cout40_9,cout40_10,cout40_11,cout40_12,cout40_13,cout41_0,cout41_1,cout41_2,cout41_3,cout41_4,cout41_5,cout41_6,cout41_7,cout41_8,cout41_9,cout41_10,cout41_11,cout41_12,cout41_13,cout42_0,cout42_1,cout42_2,cout42_3,cout42_4,cout42_5,cout42_6,cout42_7,cout42_8,cout42_9,cout42_10,cout42_11,cout42_12,cout42_13,cout43_0,cout43_1,cout43_2,cout43_3,cout43_4,cout43_5,cout43_6,cout43_7,cout43_8,cout43_9,cout43_10,cout43_11,cout43_12,cout43_13,cout44_0,cout44_1,cout44_2,cout44_3,cout44_4,cout44_5,cout44_6,cout44_7,cout44_8,cout44_9,cout44_10,cout44_11,cout44_12,cout44_13,cout45_0,cout45_1,cout45_2,cout45_3,cout45_4,cout45_5,cout45_6,cout45_7,cout45_8,cout45_9,cout45_10,cout45_11,cout45_12,cout45_13,cout46_0,cout46_1,cout46_2,cout46_3,cout46_4,cout46_5,cout46_6,cout46_7,cout46_8,cout46_9,cout46_10,cout46_11,cout46_12,cout46_13,cout47_0,cout47_1,cout47_2,cout47_3,cout47_4,cout47_5,cout47_6,cout47_7,cout47_8,cout47_9,cout47_10,cout47_11,cout47_12,cout47_13,cout48_0,cout48_1,cout48_2,cout48_3,cout48_4,cout48_5,cout48_6,cout48_7,cout48_8,cout48_9,cout48_10,cout48_11,cout48_12,cout48_13,cout49_0,cout49_1,cout49_2,cout49_3,cout49_4,cout49_5,cout49_6,cout49_7,cout49_8,cout49_9,cout49_10,cout49_11,cout49_12,cout49_13,cout50_0,cout50_1,cout50_2,cout50_3,cout50_4,cout50_5,cout50_6,cout50_7,cout50_8,cout50_9,cout50_10,cout50_11,cout50_12,cout50_13,cout51_0,cout51_1,cout51_2,cout51_3,cout51_4,cout51_5,cout51_6,cout51_7,cout51_8,cout51_9,cout51_10,cout51_11,cout51_12,cout51_13,cout52_0,cout52_1,cout52_2,cout52_3,cout52_4,cout52_5,cout52_6,cout52_7,cout52_8,cout52_9,cout52_10,cout52_11,cout52_12,cout52_13,cout53_0,cout53_1,cout53_2,cout53_3,cout53_4,cout53_5,cout53_6,cout53_7,cout53_8,cout53_9,cout53_10,cout53_11,cout53_12,cout53_13,cout54_0,cout54_1,cout54_2,cout54_3,cout54_4,cout54_5,cout54_6,cout54_7,cout54_8,cout54_9,cout54_10,cout54_11,cout54_12,cout54_13,cout55_0,cout55_1,cout55_2,cout55_3,cout55_4,cout55_5,cout55_6,cout55_7,cout55_8,cout55_9,cout55_10,cout55_11,cout55_12,cout55_13,cout56_0,cout56_1,cout56_2,cout56_3,cout56_4,cout56_5,cout56_6,cout56_7,cout56_8,cout56_9,cout56_10,cout56_11,cout56_12,cout56_13,cout57_0,cout57_1,cout57_2,cout57_3,cout57_4,cout57_5,cout57_6,cout57_7,cout57_8,cout57_9,cout57_10,cout57_11,cout57_12,cout57_13,cout58_0,cout58_1,cout58_2,cout58_3,cout58_4,cout58_5,cout58_6,cout58_7,cout58_8,cout58_9,cout58_10,cout58_11,cout58_12,cout58_13,cout59_0,cout59_1,cout59_2,cout59_3,cout59_4,cout59_5,cout59_6,cout59_7,cout59_8,cout59_9,cout59_10,cout59_11,cout59_12,cout59_13,cout60_0,cout60_1,cout60_2,cout60_3,cout60_4,cout60_5,cout60_6,cout60_7,cout60_8,cout60_9,cout60_10,cout60_11,cout60_12,cout60_13,cout61_0,cout61_1,cout61_2,cout61_3,cout61_4,cout61_5,cout61_6,cout61_7,cout61_8,cout61_9,cout61_10,cout61_11,cout61_12,cout61_13,cout62_0,cout62_1,cout62_2,cout62_3,cout62_4,cout62_5,cout62_6,cout62_7,cout62_8,cout62_9,cout62_10,cout62_11,cout62_12,cout62_13,cout63_0,cout63_1,cout63_2,cout63_3,cout63_4,cout63_5,cout63_6,cout63_7,cout63_8,cout63_9,cout63_10,cout63_11,cout63_12,cout63_13;
wire C0,C1,C2,C3,C4,C5,C6,C7,C8,C9,C10,C11,C12,C13,C14,C15,C16,C17,C18,C19,C20,C21,C22,C23,C24,C25,C26,C27,C28,C29,C30,C31,C32,C33,C34,C35,C36,C37,C38,C39,C40,C41,C42,C43,C44,C45,C46,C47,C48,C49,C50,C51,C52,C53,C54,C55,C56,C57,C58,C59,C60,C61,C62,C63;
wire S0,S1,S2,S3,S4,S5,S6,S7,S8,S9,S10,S11,S12,S13,S14,S15,S16,S17,S18,S19,S20,S21,S22,S23,S24,S25,S26,S27,S28,S29,S30,S31,S32,S33,S34,S35,S36,S37,S38,S39,S40,S41,S42,S43,S44,S45,S46,S47,S48,S49,S50,S51,S52,S53,S54,S55,S56,S57,S58,S59,S60,S61,S62,S63;

wire [63:0] in_A;
wire [63:0] in_B;
assign in_A = {S63,S62,S61,S60,S59,S58,S57,S56,S55,S54,S53,S52,S51,S50,S49,S48,S47,S46,S45,S44,S43,S42,S41,S40,S39,S38,S37,S36,S35,S34,S33,S32,S31,S30,S29,S28,S27,S26,S25,S24,S23,S22,S21,S20,S19,S18,S17,S16,S15,S14,S13,S12,S11,S10,S9,S8,S7,S6,S5,S4,S3,S2,S1,S0};
assign in_B = {C62,C61,C60,C59,C58,C57,C56,C55,C54,C53,C52,C51,C50,C49,C48,C47,C46,C45,C44,C43,C42,C41,C40,C39,C38,C37,C36,C35,C34,C33,C32,C31,C30,C29,C28,C27,C26,C25,C24,C23,C22,C21,C20,C19,C18,C17,C16,C15,C14,C13,C12,C11,C10,C9,C8,C7,C6,C5,C4,C3,C2,C1,C0,c14};

adder64 add64(
	.cin(c15),
	.A(in_A),
	.B(in_B),
	.sum(product),
	.cout()
);

//assign product = in_A + in_B;
Wallace w0(
	.n0(p0[0]),
	.n1(p1[0]),
	.n2(p2[0]),
	.n3(p3[0]),
	.n4(p4[0]),
	.n5(p5[0]),
	.n6(p6[0]),
	.n7(p7[0]),
	.n8(p8[0]),
	.n9(p9[0]),
	.n10(p10[0]),
	.n11(p11[0]),
	.n12(p12[0]),
	.n13(p13[0]),
	.n14(p14[0]),
	.n15(p15[0]),
	.cin0(c0),
	.cin1(c1),
	.cin2(c2),
	.cin3(c3),
	.cin4(c4),
	.cin5(c5),
	.cin6(c6),
	.cin7(c7),
	.cin8(c8),
	.cin9(c9),
	.cin10(c10),
	.cin11(c11),
	.cin12(c12),
	.cin13(c13),
	.c11(cout0_0),
	.c12(cout0_1),
	.c13(cout0_2),
	.c14(cout0_3),
	.c15(cout0_4),
	.c21(cout0_5),
	.c22(cout0_6),
	.c23(cout0_7),
	.c24(cout0_8),
	.c31(cout0_9),
	.c32(cout0_10),
	.c41(cout0_11),
	.c42(cout0_12),
	.c51(cout0_13),
	.c61(C0),
	.s61(S0)
);
Wallace w1(
	.n0(p0[1]),
	.n1(p1[1]),
	.n2(p2[1]),
	.n3(p3[1]),
	.n4(p4[1]),
	.n5(p5[1]),
	.n6(p6[1]),
	.n7(p7[1]),
	.n8(p8[1]),
	.n9(p9[1]),
	.n10(p10[1]),
	.n11(p11[1]),
	.n12(p12[1]),
	.n13(p13[1]),
	.n14(p14[1]),
	.n15(p15[1]),
	.cin0(cout0_0),
	.cin1(cout0_1),
	.cin2(cout0_2),
	.cin3(cout0_3),
	.cin4(cout0_4),
	.cin5(cout0_5),
	.cin6(cout0_6),
	.cin7(cout0_7),
	.cin8(cout0_8),
	.cin9(cout0_9),
	.cin10(cout0_10),
	.cin11(cout0_11),
	.cin12(cout0_12),
	.cin13(cout0_13),
	.c11(cout1_0),
	.c12(cout1_1),
	.c13(cout1_2),
	.c14(cout1_3),
	.c15(cout1_4),
	.c21(cout1_5),
	.c22(cout1_6),
	.c23(cout1_7),
	.c24(cout1_8),
	.c31(cout1_9),
	.c32(cout1_10),
	.c41(cout1_11),
	.c42(cout1_12),
	.c51(cout1_13),
	.c61(C1),
	.s61(S1)
);
Wallace w2(
	.n0(p0[2]),
	.n1(p1[2]),
	.n2(p2[2]),
	.n3(p3[2]),
	.n4(p4[2]),
	.n5(p5[2]),
	.n6(p6[2]),
	.n7(p7[2]),
	.n8(p8[2]),
	.n9(p9[2]),
	.n10(p10[2]),
	.n11(p11[2]),
	.n12(p12[2]),
	.n13(p13[2]),
	.n14(p14[2]),
	.n15(p15[2]),
	.cin0(cout1_0),
	.cin1(cout1_1),
	.cin2(cout1_2),
	.cin3(cout1_3),
	.cin4(cout1_4),
	.cin5(cout1_5),
	.cin6(cout1_6),
	.cin7(cout1_7),
	.cin8(cout1_8),
	.cin9(cout1_9),
	.cin10(cout1_10),
	.cin11(cout1_11),
	.cin12(cout1_12),
	.cin13(cout1_13),
	.c11(cout2_0),
	.c12(cout2_1),
	.c13(cout2_2),
	.c14(cout2_3),
	.c15(cout2_4),
	.c21(cout2_5),
	.c22(cout2_6),
	.c23(cout2_7),
	.c24(cout2_8),
	.c31(cout2_9),
	.c32(cout2_10),
	.c41(cout2_11),
	.c42(cout2_12),
	.c51(cout2_13),
	.c61(C2),
	.s61(S2)
);
Wallace w3(
	.n0(p0[3]),
	.n1(p1[3]),
	.n2(p2[3]),
	.n3(p3[3]),
	.n4(p4[3]),
	.n5(p5[3]),
	.n6(p6[3]),
	.n7(p7[3]),
	.n8(p8[3]),
	.n9(p9[3]),
	.n10(p10[3]),
	.n11(p11[3]),
	.n12(p12[3]),
	.n13(p13[3]),
	.n14(p14[3]),
	.n15(p15[3]),
	.cin0(cout2_0),
	.cin1(cout2_1),
	.cin2(cout2_2),
	.cin3(cout2_3),
	.cin4(cout2_4),
	.cin5(cout2_5),
	.cin6(cout2_6),
	.cin7(cout2_7),
	.cin8(cout2_8),
	.cin9(cout2_9),
	.cin10(cout2_10),
	.cin11(cout2_11),
	.cin12(cout2_12),
	.cin13(cout2_13),
	.c11(cout3_0),
	.c12(cout3_1),
	.c13(cout3_2),
	.c14(cout3_3),
	.c15(cout3_4),
	.c21(cout3_5),
	.c22(cout3_6),
	.c23(cout3_7),
	.c24(cout3_8),
	.c31(cout3_9),
	.c32(cout3_10),
	.c41(cout3_11),
	.c42(cout3_12),
	.c51(cout3_13),
	.c61(C3),
	.s61(S3)
);
Wallace w4(
	.n0(p0[4]),
	.n1(p1[4]),
	.n2(p2[4]),
	.n3(p3[4]),
	.n4(p4[4]),
	.n5(p5[4]),
	.n6(p6[4]),
	.n7(p7[4]),
	.n8(p8[4]),
	.n9(p9[4]),
	.n10(p10[4]),
	.n11(p11[4]),
	.n12(p12[4]),
	.n13(p13[4]),
	.n14(p14[4]),
	.n15(p15[4]),
	.cin0(cout3_0),
	.cin1(cout3_1),
	.cin2(cout3_2),
	.cin3(cout3_3),
	.cin4(cout3_4),
	.cin5(cout3_5),
	.cin6(cout3_6),
	.cin7(cout3_7),
	.cin8(cout3_8),
	.cin9(cout3_9),
	.cin10(cout3_10),
	.cin11(cout3_11),
	.cin12(cout3_12),
	.cin13(cout3_13),
	.c11(cout4_0),
	.c12(cout4_1),
	.c13(cout4_2),
	.c14(cout4_3),
	.c15(cout4_4),
	.c21(cout4_5),
	.c22(cout4_6),
	.c23(cout4_7),
	.c24(cout4_8),
	.c31(cout4_9),
	.c32(cout4_10),
	.c41(cout4_11),
	.c42(cout4_12),
	.c51(cout4_13),
	.c61(C4),
	.s61(S4)
);
Wallace w5(
	.n0(p0[5]),
	.n1(p1[5]),
	.n2(p2[5]),
	.n3(p3[5]),
	.n4(p4[5]),
	.n5(p5[5]),
	.n6(p6[5]),
	.n7(p7[5]),
	.n8(p8[5]),
	.n9(p9[5]),
	.n10(p10[5]),
	.n11(p11[5]),
	.n12(p12[5]),
	.n13(p13[5]),
	.n14(p14[5]),
	.n15(p15[5]),
	.cin0(cout4_0),
	.cin1(cout4_1),
	.cin2(cout4_2),
	.cin3(cout4_3),
	.cin4(cout4_4),
	.cin5(cout4_5),
	.cin6(cout4_6),
	.cin7(cout4_7),
	.cin8(cout4_8),
	.cin9(cout4_9),
	.cin10(cout4_10),
	.cin11(cout4_11),
	.cin12(cout4_12),
	.cin13(cout4_13),
	.c11(cout5_0),
	.c12(cout5_1),
	.c13(cout5_2),
	.c14(cout5_3),
	.c15(cout5_4),
	.c21(cout5_5),
	.c22(cout5_6),
	.c23(cout5_7),
	.c24(cout5_8),
	.c31(cout5_9),
	.c32(cout5_10),
	.c41(cout5_11),
	.c42(cout5_12),
	.c51(cout5_13),
	.c61(C5),
	.s61(S5)
);
Wallace w6(
	.n0(p0[6]),
	.n1(p1[6]),
	.n2(p2[6]),
	.n3(p3[6]),
	.n4(p4[6]),
	.n5(p5[6]),
	.n6(p6[6]),
	.n7(p7[6]),
	.n8(p8[6]),
	.n9(p9[6]),
	.n10(p10[6]),
	.n11(p11[6]),
	.n12(p12[6]),
	.n13(p13[6]),
	.n14(p14[6]),
	.n15(p15[6]),
	.cin0(cout5_0),
	.cin1(cout5_1),
	.cin2(cout5_2),
	.cin3(cout5_3),
	.cin4(cout5_4),
	.cin5(cout5_5),
	.cin6(cout5_6),
	.cin7(cout5_7),
	.cin8(cout5_8),
	.cin9(cout5_9),
	.cin10(cout5_10),
	.cin11(cout5_11),
	.cin12(cout5_12),
	.cin13(cout5_13),
	.c11(cout6_0),
	.c12(cout6_1),
	.c13(cout6_2),
	.c14(cout6_3),
	.c15(cout6_4),
	.c21(cout6_5),
	.c22(cout6_6),
	.c23(cout6_7),
	.c24(cout6_8),
	.c31(cout6_9),
	.c32(cout6_10),
	.c41(cout6_11),
	.c42(cout6_12),
	.c51(cout6_13),
	.c61(C6),
	.s61(S6)
);
Wallace w7(
	.n0(p0[7]),
	.n1(p1[7]),
	.n2(p2[7]),
	.n3(p3[7]),
	.n4(p4[7]),
	.n5(p5[7]),
	.n6(p6[7]),
	.n7(p7[7]),
	.n8(p8[7]),
	.n9(p9[7]),
	.n10(p10[7]),
	.n11(p11[7]),
	.n12(p12[7]),
	.n13(p13[7]),
	.n14(p14[7]),
	.n15(p15[7]),
	.cin0(cout6_0),
	.cin1(cout6_1),
	.cin2(cout6_2),
	.cin3(cout6_3),
	.cin4(cout6_4),
	.cin5(cout6_5),
	.cin6(cout6_6),
	.cin7(cout6_7),
	.cin8(cout6_8),
	.cin9(cout6_9),
	.cin10(cout6_10),
	.cin11(cout6_11),
	.cin12(cout6_12),
	.cin13(cout6_13),
	.c11(cout7_0),
	.c12(cout7_1),
	.c13(cout7_2),
	.c14(cout7_3),
	.c15(cout7_4),
	.c21(cout7_5),
	.c22(cout7_6),
	.c23(cout7_7),
	.c24(cout7_8),
	.c31(cout7_9),
	.c32(cout7_10),
	.c41(cout7_11),
	.c42(cout7_12),
	.c51(cout7_13),
	.c61(C7),
	.s61(S7)
);
Wallace w8(
	.n0(p0[8]),
	.n1(p1[8]),
	.n2(p2[8]),
	.n3(p3[8]),
	.n4(p4[8]),
	.n5(p5[8]),
	.n6(p6[8]),
	.n7(p7[8]),
	.n8(p8[8]),
	.n9(p9[8]),
	.n10(p10[8]),
	.n11(p11[8]),
	.n12(p12[8]),
	.n13(p13[8]),
	.n14(p14[8]),
	.n15(p15[8]),
	.cin0(cout7_0),
	.cin1(cout7_1),
	.cin2(cout7_2),
	.cin3(cout7_3),
	.cin4(cout7_4),
	.cin5(cout7_5),
	.cin6(cout7_6),
	.cin7(cout7_7),
	.cin8(cout7_8),
	.cin9(cout7_9),
	.cin10(cout7_10),
	.cin11(cout7_11),
	.cin12(cout7_12),
	.cin13(cout7_13),
	.c11(cout8_0),
	.c12(cout8_1),
	.c13(cout8_2),
	.c14(cout8_3),
	.c15(cout8_4),
	.c21(cout8_5),
	.c22(cout8_6),
	.c23(cout8_7),
	.c24(cout8_8),
	.c31(cout8_9),
	.c32(cout8_10),
	.c41(cout8_11),
	.c42(cout8_12),
	.c51(cout8_13),
	.c61(C8),
	.s61(S8)
);
Wallace w9(
	.n0(p0[9]),
	.n1(p1[9]),
	.n2(p2[9]),
	.n3(p3[9]),
	.n4(p4[9]),
	.n5(p5[9]),
	.n6(p6[9]),
	.n7(p7[9]),
	.n8(p8[9]),
	.n9(p9[9]),
	.n10(p10[9]),
	.n11(p11[9]),
	.n12(p12[9]),
	.n13(p13[9]),
	.n14(p14[9]),
	.n15(p15[9]),
	.cin0(cout8_0),
	.cin1(cout8_1),
	.cin2(cout8_2),
	.cin3(cout8_3),
	.cin4(cout8_4),
	.cin5(cout8_5),
	.cin6(cout8_6),
	.cin7(cout8_7),
	.cin8(cout8_8),
	.cin9(cout8_9),
	.cin10(cout8_10),
	.cin11(cout8_11),
	.cin12(cout8_12),
	.cin13(cout8_13),
	.c11(cout9_0),
	.c12(cout9_1),
	.c13(cout9_2),
	.c14(cout9_3),
	.c15(cout9_4),
	.c21(cout9_5),
	.c22(cout9_6),
	.c23(cout9_7),
	.c24(cout9_8),
	.c31(cout9_9),
	.c32(cout9_10),
	.c41(cout9_11),
	.c42(cout9_12),
	.c51(cout9_13),
	.c61(C9),
	.s61(S9)
);
Wallace w10(
	.n0(p0[10]),
	.n1(p1[10]),
	.n2(p2[10]),
	.n3(p3[10]),
	.n4(p4[10]),
	.n5(p5[10]),
	.n6(p6[10]),
	.n7(p7[10]),
	.n8(p8[10]),
	.n9(p9[10]),
	.n10(p10[10]),
	.n11(p11[10]),
	.n12(p12[10]),
	.n13(p13[10]),
	.n14(p14[10]),
	.n15(p15[10]),
	.cin0(cout9_0),
	.cin1(cout9_1),
	.cin2(cout9_2),
	.cin3(cout9_3),
	.cin4(cout9_4),
	.cin5(cout9_5),
	.cin6(cout9_6),
	.cin7(cout9_7),
	.cin8(cout9_8),
	.cin9(cout9_9),
	.cin10(cout9_10),
	.cin11(cout9_11),
	.cin12(cout9_12),
	.cin13(cout9_13),
	.c11(cout10_0),
	.c12(cout10_1),
	.c13(cout10_2),
	.c14(cout10_3),
	.c15(cout10_4),
	.c21(cout10_5),
	.c22(cout10_6),
	.c23(cout10_7),
	.c24(cout10_8),
	.c31(cout10_9),
	.c32(cout10_10),
	.c41(cout10_11),
	.c42(cout10_12),
	.c51(cout10_13),
	.c61(C10),
	.s61(S10)
);
Wallace w11(
	.n0(p0[11]),
	.n1(p1[11]),
	.n2(p2[11]),
	.n3(p3[11]),
	.n4(p4[11]),
	.n5(p5[11]),
	.n6(p6[11]),
	.n7(p7[11]),
	.n8(p8[11]),
	.n9(p9[11]),
	.n10(p10[11]),
	.n11(p11[11]),
	.n12(p12[11]),
	.n13(p13[11]),
	.n14(p14[11]),
	.n15(p15[11]),
	.cin0(cout10_0),
	.cin1(cout10_1),
	.cin2(cout10_2),
	.cin3(cout10_3),
	.cin4(cout10_4),
	.cin5(cout10_5),
	.cin6(cout10_6),
	.cin7(cout10_7),
	.cin8(cout10_8),
	.cin9(cout10_9),
	.cin10(cout10_10),
	.cin11(cout10_11),
	.cin12(cout10_12),
	.cin13(cout10_13),
	.c11(cout11_0),
	.c12(cout11_1),
	.c13(cout11_2),
	.c14(cout11_3),
	.c15(cout11_4),
	.c21(cout11_5),
	.c22(cout11_6),
	.c23(cout11_7),
	.c24(cout11_8),
	.c31(cout11_9),
	.c32(cout11_10),
	.c41(cout11_11),
	.c42(cout11_12),
	.c51(cout11_13),
	.c61(C11),
	.s61(S11)
);
Wallace w12(
	.n0(p0[12]),
	.n1(p1[12]),
	.n2(p2[12]),
	.n3(p3[12]),
	.n4(p4[12]),
	.n5(p5[12]),
	.n6(p6[12]),
	.n7(p7[12]),
	.n8(p8[12]),
	.n9(p9[12]),
	.n10(p10[12]),
	.n11(p11[12]),
	.n12(p12[12]),
	.n13(p13[12]),
	.n14(p14[12]),
	.n15(p15[12]),
	.cin0(cout11_0),
	.cin1(cout11_1),
	.cin2(cout11_2),
	.cin3(cout11_3),
	.cin4(cout11_4),
	.cin5(cout11_5),
	.cin6(cout11_6),
	.cin7(cout11_7),
	.cin8(cout11_8),
	.cin9(cout11_9),
	.cin10(cout11_10),
	.cin11(cout11_11),
	.cin12(cout11_12),
	.cin13(cout11_13),
	.c11(cout12_0),
	.c12(cout12_1),
	.c13(cout12_2),
	.c14(cout12_3),
	.c15(cout12_4),
	.c21(cout12_5),
	.c22(cout12_6),
	.c23(cout12_7),
	.c24(cout12_8),
	.c31(cout12_9),
	.c32(cout12_10),
	.c41(cout12_11),
	.c42(cout12_12),
	.c51(cout12_13),
	.c61(C12),
	.s61(S12)
);
Wallace w13(
	.n0(p0[13]),
	.n1(p1[13]),
	.n2(p2[13]),
	.n3(p3[13]),
	.n4(p4[13]),
	.n5(p5[13]),
	.n6(p6[13]),
	.n7(p7[13]),
	.n8(p8[13]),
	.n9(p9[13]),
	.n10(p10[13]),
	.n11(p11[13]),
	.n12(p12[13]),
	.n13(p13[13]),
	.n14(p14[13]),
	.n15(p15[13]),
	.cin0(cout12_0),
	.cin1(cout12_1),
	.cin2(cout12_2),
	.cin3(cout12_3),
	.cin4(cout12_4),
	.cin5(cout12_5),
	.cin6(cout12_6),
	.cin7(cout12_7),
	.cin8(cout12_8),
	.cin9(cout12_9),
	.cin10(cout12_10),
	.cin11(cout12_11),
	.cin12(cout12_12),
	.cin13(cout12_13),
	.c11(cout13_0),
	.c12(cout13_1),
	.c13(cout13_2),
	.c14(cout13_3),
	.c15(cout13_4),
	.c21(cout13_5),
	.c22(cout13_6),
	.c23(cout13_7),
	.c24(cout13_8),
	.c31(cout13_9),
	.c32(cout13_10),
	.c41(cout13_11),
	.c42(cout13_12),
	.c51(cout13_13),
	.c61(C13),
	.s61(S13)
);
Wallace w14(
	.n0(p0[14]),
	.n1(p1[14]),
	.n2(p2[14]),
	.n3(p3[14]),
	.n4(p4[14]),
	.n5(p5[14]),
	.n6(p6[14]),
	.n7(p7[14]),
	.n8(p8[14]),
	.n9(p9[14]),
	.n10(p10[14]),
	.n11(p11[14]),
	.n12(p12[14]),
	.n13(p13[14]),
	.n14(p14[14]),
	.n15(p15[14]),
	.cin0(cout13_0),
	.cin1(cout13_1),
	.cin2(cout13_2),
	.cin3(cout13_3),
	.cin4(cout13_4),
	.cin5(cout13_5),
	.cin6(cout13_6),
	.cin7(cout13_7),
	.cin8(cout13_8),
	.cin9(cout13_9),
	.cin10(cout13_10),
	.cin11(cout13_11),
	.cin12(cout13_12),
	.cin13(cout13_13),
	.c11(cout14_0),
	.c12(cout14_1),
	.c13(cout14_2),
	.c14(cout14_3),
	.c15(cout14_4),
	.c21(cout14_5),
	.c22(cout14_6),
	.c23(cout14_7),
	.c24(cout14_8),
	.c31(cout14_9),
	.c32(cout14_10),
	.c41(cout14_11),
	.c42(cout14_12),
	.c51(cout14_13),
	.c61(C14),
	.s61(S14)
);
Wallace w15(
	.n0(p0[15]),
	.n1(p1[15]),
	.n2(p2[15]),
	.n3(p3[15]),
	.n4(p4[15]),
	.n5(p5[15]),
	.n6(p6[15]),
	.n7(p7[15]),
	.n8(p8[15]),
	.n9(p9[15]),
	.n10(p10[15]),
	.n11(p11[15]),
	.n12(p12[15]),
	.n13(p13[15]),
	.n14(p14[15]),
	.n15(p15[15]),
	.cin0(cout14_0),
	.cin1(cout14_1),
	.cin2(cout14_2),
	.cin3(cout14_3),
	.cin4(cout14_4),
	.cin5(cout14_5),
	.cin6(cout14_6),
	.cin7(cout14_7),
	.cin8(cout14_8),
	.cin9(cout14_9),
	.cin10(cout14_10),
	.cin11(cout14_11),
	.cin12(cout14_12),
	.cin13(cout14_13),
	.c11(cout15_0),
	.c12(cout15_1),
	.c13(cout15_2),
	.c14(cout15_3),
	.c15(cout15_4),
	.c21(cout15_5),
	.c22(cout15_6),
	.c23(cout15_7),
	.c24(cout15_8),
	.c31(cout15_9),
	.c32(cout15_10),
	.c41(cout15_11),
	.c42(cout15_12),
	.c51(cout15_13),
	.c61(C15),
	.s61(S15)
);
Wallace w16(
	.n0(p0[16]),
	.n1(p1[16]),
	.n2(p2[16]),
	.n3(p3[16]),
	.n4(p4[16]),
	.n5(p5[16]),
	.n6(p6[16]),
	.n7(p7[16]),
	.n8(p8[16]),
	.n9(p9[16]),
	.n10(p10[16]),
	.n11(p11[16]),
	.n12(p12[16]),
	.n13(p13[16]),
	.n14(p14[16]),
	.n15(p15[16]),
	.cin0(cout15_0),
	.cin1(cout15_1),
	.cin2(cout15_2),
	.cin3(cout15_3),
	.cin4(cout15_4),
	.cin5(cout15_5),
	.cin6(cout15_6),
	.cin7(cout15_7),
	.cin8(cout15_8),
	.cin9(cout15_9),
	.cin10(cout15_10),
	.cin11(cout15_11),
	.cin12(cout15_12),
	.cin13(cout15_13),
	.c11(cout16_0),
	.c12(cout16_1),
	.c13(cout16_2),
	.c14(cout16_3),
	.c15(cout16_4),
	.c21(cout16_5),
	.c22(cout16_6),
	.c23(cout16_7),
	.c24(cout16_8),
	.c31(cout16_9),
	.c32(cout16_10),
	.c41(cout16_11),
	.c42(cout16_12),
	.c51(cout16_13),
	.c61(C16),
	.s61(S16)
);
Wallace w17(
	.n0(p0[17]),
	.n1(p1[17]),
	.n2(p2[17]),
	.n3(p3[17]),
	.n4(p4[17]),
	.n5(p5[17]),
	.n6(p6[17]),
	.n7(p7[17]),
	.n8(p8[17]),
	.n9(p9[17]),
	.n10(p10[17]),
	.n11(p11[17]),
	.n12(p12[17]),
	.n13(p13[17]),
	.n14(p14[17]),
	.n15(p15[17]),
	.cin0(cout16_0),
	.cin1(cout16_1),
	.cin2(cout16_2),
	.cin3(cout16_3),
	.cin4(cout16_4),
	.cin5(cout16_5),
	.cin6(cout16_6),
	.cin7(cout16_7),
	.cin8(cout16_8),
	.cin9(cout16_9),
	.cin10(cout16_10),
	.cin11(cout16_11),
	.cin12(cout16_12),
	.cin13(cout16_13),
	.c11(cout17_0),
	.c12(cout17_1),
	.c13(cout17_2),
	.c14(cout17_3),
	.c15(cout17_4),
	.c21(cout17_5),
	.c22(cout17_6),
	.c23(cout17_7),
	.c24(cout17_8),
	.c31(cout17_9),
	.c32(cout17_10),
	.c41(cout17_11),
	.c42(cout17_12),
	.c51(cout17_13),
	.c61(C17),
	.s61(S17)
);
Wallace w18(
	.n0(p0[18]),
	.n1(p1[18]),
	.n2(p2[18]),
	.n3(p3[18]),
	.n4(p4[18]),
	.n5(p5[18]),
	.n6(p6[18]),
	.n7(p7[18]),
	.n8(p8[18]),
	.n9(p9[18]),
	.n10(p10[18]),
	.n11(p11[18]),
	.n12(p12[18]),
	.n13(p13[18]),
	.n14(p14[18]),
	.n15(p15[18]),
	.cin0(cout17_0),
	.cin1(cout17_1),
	.cin2(cout17_2),
	.cin3(cout17_3),
	.cin4(cout17_4),
	.cin5(cout17_5),
	.cin6(cout17_6),
	.cin7(cout17_7),
	.cin8(cout17_8),
	.cin9(cout17_9),
	.cin10(cout17_10),
	.cin11(cout17_11),
	.cin12(cout17_12),
	.cin13(cout17_13),
	.c11(cout18_0),
	.c12(cout18_1),
	.c13(cout18_2),
	.c14(cout18_3),
	.c15(cout18_4),
	.c21(cout18_5),
	.c22(cout18_6),
	.c23(cout18_7),
	.c24(cout18_8),
	.c31(cout18_9),
	.c32(cout18_10),
	.c41(cout18_11),
	.c42(cout18_12),
	.c51(cout18_13),
	.c61(C18),
	.s61(S18)
);
Wallace w19(
	.n0(p0[19]),
	.n1(p1[19]),
	.n2(p2[19]),
	.n3(p3[19]),
	.n4(p4[19]),
	.n5(p5[19]),
	.n6(p6[19]),
	.n7(p7[19]),
	.n8(p8[19]),
	.n9(p9[19]),
	.n10(p10[19]),
	.n11(p11[19]),
	.n12(p12[19]),
	.n13(p13[19]),
	.n14(p14[19]),
	.n15(p15[19]),
	.cin0(cout18_0),
	.cin1(cout18_1),
	.cin2(cout18_2),
	.cin3(cout18_3),
	.cin4(cout18_4),
	.cin5(cout18_5),
	.cin6(cout18_6),
	.cin7(cout18_7),
	.cin8(cout18_8),
	.cin9(cout18_9),
	.cin10(cout18_10),
	.cin11(cout18_11),
	.cin12(cout18_12),
	.cin13(cout18_13),
	.c11(cout19_0),
	.c12(cout19_1),
	.c13(cout19_2),
	.c14(cout19_3),
	.c15(cout19_4),
	.c21(cout19_5),
	.c22(cout19_6),
	.c23(cout19_7),
	.c24(cout19_8),
	.c31(cout19_9),
	.c32(cout19_10),
	.c41(cout19_11),
	.c42(cout19_12),
	.c51(cout19_13),
	.c61(C19),
	.s61(S19)
);
Wallace w20(
	.n0(p0[20]),
	.n1(p1[20]),
	.n2(p2[20]),
	.n3(p3[20]),
	.n4(p4[20]),
	.n5(p5[20]),
	.n6(p6[20]),
	.n7(p7[20]),
	.n8(p8[20]),
	.n9(p9[20]),
	.n10(p10[20]),
	.n11(p11[20]),
	.n12(p12[20]),
	.n13(p13[20]),
	.n14(p14[20]),
	.n15(p15[20]),
	.cin0(cout19_0),
	.cin1(cout19_1),
	.cin2(cout19_2),
	.cin3(cout19_3),
	.cin4(cout19_4),
	.cin5(cout19_5),
	.cin6(cout19_6),
	.cin7(cout19_7),
	.cin8(cout19_8),
	.cin9(cout19_9),
	.cin10(cout19_10),
	.cin11(cout19_11),
	.cin12(cout19_12),
	.cin13(cout19_13),
	.c11(cout20_0),
	.c12(cout20_1),
	.c13(cout20_2),
	.c14(cout20_3),
	.c15(cout20_4),
	.c21(cout20_5),
	.c22(cout20_6),
	.c23(cout20_7),
	.c24(cout20_8),
	.c31(cout20_9),
	.c32(cout20_10),
	.c41(cout20_11),
	.c42(cout20_12),
	.c51(cout20_13),
	.c61(C20),
	.s61(S20)
);
Wallace w21(
	.n0(p0[21]),
	.n1(p1[21]),
	.n2(p2[21]),
	.n3(p3[21]),
	.n4(p4[21]),
	.n5(p5[21]),
	.n6(p6[21]),
	.n7(p7[21]),
	.n8(p8[21]),
	.n9(p9[21]),
	.n10(p10[21]),
	.n11(p11[21]),
	.n12(p12[21]),
	.n13(p13[21]),
	.n14(p14[21]),
	.n15(p15[21]),
	.cin0(cout20_0),
	.cin1(cout20_1),
	.cin2(cout20_2),
	.cin3(cout20_3),
	.cin4(cout20_4),
	.cin5(cout20_5),
	.cin6(cout20_6),
	.cin7(cout20_7),
	.cin8(cout20_8),
	.cin9(cout20_9),
	.cin10(cout20_10),
	.cin11(cout20_11),
	.cin12(cout20_12),
	.cin13(cout20_13),
	.c11(cout21_0),
	.c12(cout21_1),
	.c13(cout21_2),
	.c14(cout21_3),
	.c15(cout21_4),
	.c21(cout21_5),
	.c22(cout21_6),
	.c23(cout21_7),
	.c24(cout21_8),
	.c31(cout21_9),
	.c32(cout21_10),
	.c41(cout21_11),
	.c42(cout21_12),
	.c51(cout21_13),
	.c61(C21),
	.s61(S21)
);
Wallace w22(
	.n0(p0[22]),
	.n1(p1[22]),
	.n2(p2[22]),
	.n3(p3[22]),
	.n4(p4[22]),
	.n5(p5[22]),
	.n6(p6[22]),
	.n7(p7[22]),
	.n8(p8[22]),
	.n9(p9[22]),
	.n10(p10[22]),
	.n11(p11[22]),
	.n12(p12[22]),
	.n13(p13[22]),
	.n14(p14[22]),
	.n15(p15[22]),
	.cin0(cout21_0),
	.cin1(cout21_1),
	.cin2(cout21_2),
	.cin3(cout21_3),
	.cin4(cout21_4),
	.cin5(cout21_5),
	.cin6(cout21_6),
	.cin7(cout21_7),
	.cin8(cout21_8),
	.cin9(cout21_9),
	.cin10(cout21_10),
	.cin11(cout21_11),
	.cin12(cout21_12),
	.cin13(cout21_13),
	.c11(cout22_0),
	.c12(cout22_1),
	.c13(cout22_2),
	.c14(cout22_3),
	.c15(cout22_4),
	.c21(cout22_5),
	.c22(cout22_6),
	.c23(cout22_7),
	.c24(cout22_8),
	.c31(cout22_9),
	.c32(cout22_10),
	.c41(cout22_11),
	.c42(cout22_12),
	.c51(cout22_13),
	.c61(C22),
	.s61(S22)
);
Wallace w23(
	.n0(p0[23]),
	.n1(p1[23]),
	.n2(p2[23]),
	.n3(p3[23]),
	.n4(p4[23]),
	.n5(p5[23]),
	.n6(p6[23]),
	.n7(p7[23]),
	.n8(p8[23]),
	.n9(p9[23]),
	.n10(p10[23]),
	.n11(p11[23]),
	.n12(p12[23]),
	.n13(p13[23]),
	.n14(p14[23]),
	.n15(p15[23]),
	.cin0(cout22_0),
	.cin1(cout22_1),
	.cin2(cout22_2),
	.cin3(cout22_3),
	.cin4(cout22_4),
	.cin5(cout22_5),
	.cin6(cout22_6),
	.cin7(cout22_7),
	.cin8(cout22_8),
	.cin9(cout22_9),
	.cin10(cout22_10),
	.cin11(cout22_11),
	.cin12(cout22_12),
	.cin13(cout22_13),
	.c11(cout23_0),
	.c12(cout23_1),
	.c13(cout23_2),
	.c14(cout23_3),
	.c15(cout23_4),
	.c21(cout23_5),
	.c22(cout23_6),
	.c23(cout23_7),
	.c24(cout23_8),
	.c31(cout23_9),
	.c32(cout23_10),
	.c41(cout23_11),
	.c42(cout23_12),
	.c51(cout23_13),
	.c61(C23),
	.s61(S23)
);
Wallace w24(
	.n0(p0[24]),
	.n1(p1[24]),
	.n2(p2[24]),
	.n3(p3[24]),
	.n4(p4[24]),
	.n5(p5[24]),
	.n6(p6[24]),
	.n7(p7[24]),
	.n8(p8[24]),
	.n9(p9[24]),
	.n10(p10[24]),
	.n11(p11[24]),
	.n12(p12[24]),
	.n13(p13[24]),
	.n14(p14[24]),
	.n15(p15[24]),
	.cin0(cout23_0),
	.cin1(cout23_1),
	.cin2(cout23_2),
	.cin3(cout23_3),
	.cin4(cout23_4),
	.cin5(cout23_5),
	.cin6(cout23_6),
	.cin7(cout23_7),
	.cin8(cout23_8),
	.cin9(cout23_9),
	.cin10(cout23_10),
	.cin11(cout23_11),
	.cin12(cout23_12),
	.cin13(cout23_13),
	.c11(cout24_0),
	.c12(cout24_1),
	.c13(cout24_2),
	.c14(cout24_3),
	.c15(cout24_4),
	.c21(cout24_5),
	.c22(cout24_6),
	.c23(cout24_7),
	.c24(cout24_8),
	.c31(cout24_9),
	.c32(cout24_10),
	.c41(cout24_11),
	.c42(cout24_12),
	.c51(cout24_13),
	.c61(C24),
	.s61(S24)
);
Wallace w25(
	.n0(p0[25]),
	.n1(p1[25]),
	.n2(p2[25]),
	.n3(p3[25]),
	.n4(p4[25]),
	.n5(p5[25]),
	.n6(p6[25]),
	.n7(p7[25]),
	.n8(p8[25]),
	.n9(p9[25]),
	.n10(p10[25]),
	.n11(p11[25]),
	.n12(p12[25]),
	.n13(p13[25]),
	.n14(p14[25]),
	.n15(p15[25]),
	.cin0(cout24_0),
	.cin1(cout24_1),
	.cin2(cout24_2),
	.cin3(cout24_3),
	.cin4(cout24_4),
	.cin5(cout24_5),
	.cin6(cout24_6),
	.cin7(cout24_7),
	.cin8(cout24_8),
	.cin9(cout24_9),
	.cin10(cout24_10),
	.cin11(cout24_11),
	.cin12(cout24_12),
	.cin13(cout24_13),
	.c11(cout25_0),
	.c12(cout25_1),
	.c13(cout25_2),
	.c14(cout25_3),
	.c15(cout25_4),
	.c21(cout25_5),
	.c22(cout25_6),
	.c23(cout25_7),
	.c24(cout25_8),
	.c31(cout25_9),
	.c32(cout25_10),
	.c41(cout25_11),
	.c42(cout25_12),
	.c51(cout25_13),
	.c61(C25),
	.s61(S25)
);
Wallace w26(
	.n0(p0[26]),
	.n1(p1[26]),
	.n2(p2[26]),
	.n3(p3[26]),
	.n4(p4[26]),
	.n5(p5[26]),
	.n6(p6[26]),
	.n7(p7[26]),
	.n8(p8[26]),
	.n9(p9[26]),
	.n10(p10[26]),
	.n11(p11[26]),
	.n12(p12[26]),
	.n13(p13[26]),
	.n14(p14[26]),
	.n15(p15[26]),
	.cin0(cout25_0),
	.cin1(cout25_1),
	.cin2(cout25_2),
	.cin3(cout25_3),
	.cin4(cout25_4),
	.cin5(cout25_5),
	.cin6(cout25_6),
	.cin7(cout25_7),
	.cin8(cout25_8),
	.cin9(cout25_9),
	.cin10(cout25_10),
	.cin11(cout25_11),
	.cin12(cout25_12),
	.cin13(cout25_13),
	.c11(cout26_0),
	.c12(cout26_1),
	.c13(cout26_2),
	.c14(cout26_3),
	.c15(cout26_4),
	.c21(cout26_5),
	.c22(cout26_6),
	.c23(cout26_7),
	.c24(cout26_8),
	.c31(cout26_9),
	.c32(cout26_10),
	.c41(cout26_11),
	.c42(cout26_12),
	.c51(cout26_13),
	.c61(C26),
	.s61(S26)
);
Wallace w27(
	.n0(p0[27]),
	.n1(p1[27]),
	.n2(p2[27]),
	.n3(p3[27]),
	.n4(p4[27]),
	.n5(p5[27]),
	.n6(p6[27]),
	.n7(p7[27]),
	.n8(p8[27]),
	.n9(p9[27]),
	.n10(p10[27]),
	.n11(p11[27]),
	.n12(p12[27]),
	.n13(p13[27]),
	.n14(p14[27]),
	.n15(p15[27]),
	.cin0(cout26_0),
	.cin1(cout26_1),
	.cin2(cout26_2),
	.cin3(cout26_3),
	.cin4(cout26_4),
	.cin5(cout26_5),
	.cin6(cout26_6),
	.cin7(cout26_7),
	.cin8(cout26_8),
	.cin9(cout26_9),
	.cin10(cout26_10),
	.cin11(cout26_11),
	.cin12(cout26_12),
	.cin13(cout26_13),
	.c11(cout27_0),
	.c12(cout27_1),
	.c13(cout27_2),
	.c14(cout27_3),
	.c15(cout27_4),
	.c21(cout27_5),
	.c22(cout27_6),
	.c23(cout27_7),
	.c24(cout27_8),
	.c31(cout27_9),
	.c32(cout27_10),
	.c41(cout27_11),
	.c42(cout27_12),
	.c51(cout27_13),
	.c61(C27),
	.s61(S27)
);
Wallace w28(
	.n0(p0[28]),
	.n1(p1[28]),
	.n2(p2[28]),
	.n3(p3[28]),
	.n4(p4[28]),
	.n5(p5[28]),
	.n6(p6[28]),
	.n7(p7[28]),
	.n8(p8[28]),
	.n9(p9[28]),
	.n10(p10[28]),
	.n11(p11[28]),
	.n12(p12[28]),
	.n13(p13[28]),
	.n14(p14[28]),
	.n15(p15[28]),
	.cin0(cout27_0),
	.cin1(cout27_1),
	.cin2(cout27_2),
	.cin3(cout27_3),
	.cin4(cout27_4),
	.cin5(cout27_5),
	.cin6(cout27_6),
	.cin7(cout27_7),
	.cin8(cout27_8),
	.cin9(cout27_9),
	.cin10(cout27_10),
	.cin11(cout27_11),
	.cin12(cout27_12),
	.cin13(cout27_13),
	.c11(cout28_0),
	.c12(cout28_1),
	.c13(cout28_2),
	.c14(cout28_3),
	.c15(cout28_4),
	.c21(cout28_5),
	.c22(cout28_6),
	.c23(cout28_7),
	.c24(cout28_8),
	.c31(cout28_9),
	.c32(cout28_10),
	.c41(cout28_11),
	.c42(cout28_12),
	.c51(cout28_13),
	.c61(C28),
	.s61(S28)
);
Wallace w29(
	.n0(p0[29]),
	.n1(p1[29]),
	.n2(p2[29]),
	.n3(p3[29]),
	.n4(p4[29]),
	.n5(p5[29]),
	.n6(p6[29]),
	.n7(p7[29]),
	.n8(p8[29]),
	.n9(p9[29]),
	.n10(p10[29]),
	.n11(p11[29]),
	.n12(p12[29]),
	.n13(p13[29]),
	.n14(p14[29]),
	.n15(p15[29]),
	.cin0(cout28_0),
	.cin1(cout28_1),
	.cin2(cout28_2),
	.cin3(cout28_3),
	.cin4(cout28_4),
	.cin5(cout28_5),
	.cin6(cout28_6),
	.cin7(cout28_7),
	.cin8(cout28_8),
	.cin9(cout28_9),
	.cin10(cout28_10),
	.cin11(cout28_11),
	.cin12(cout28_12),
	.cin13(cout28_13),
	.c11(cout29_0),
	.c12(cout29_1),
	.c13(cout29_2),
	.c14(cout29_3),
	.c15(cout29_4),
	.c21(cout29_5),
	.c22(cout29_6),
	.c23(cout29_7),
	.c24(cout29_8),
	.c31(cout29_9),
	.c32(cout29_10),
	.c41(cout29_11),
	.c42(cout29_12),
	.c51(cout29_13),
	.c61(C29),
	.s61(S29)
);
Wallace w30(
	.n0(p0[30]),
	.n1(p1[30]),
	.n2(p2[30]),
	.n3(p3[30]),
	.n4(p4[30]),
	.n5(p5[30]),
	.n6(p6[30]),
	.n7(p7[30]),
	.n8(p8[30]),
	.n9(p9[30]),
	.n10(p10[30]),
	.n11(p11[30]),
	.n12(p12[30]),
	.n13(p13[30]),
	.n14(p14[30]),
	.n15(p15[30]),
	.cin0(cout29_0),
	.cin1(cout29_1),
	.cin2(cout29_2),
	.cin3(cout29_3),
	.cin4(cout29_4),
	.cin5(cout29_5),
	.cin6(cout29_6),
	.cin7(cout29_7),
	.cin8(cout29_8),
	.cin9(cout29_9),
	.cin10(cout29_10),
	.cin11(cout29_11),
	.cin12(cout29_12),
	.cin13(cout29_13),
	.c11(cout30_0),
	.c12(cout30_1),
	.c13(cout30_2),
	.c14(cout30_3),
	.c15(cout30_4),
	.c21(cout30_5),
	.c22(cout30_6),
	.c23(cout30_7),
	.c24(cout30_8),
	.c31(cout30_9),
	.c32(cout30_10),
	.c41(cout30_11),
	.c42(cout30_12),
	.c51(cout30_13),
	.c61(C30),
	.s61(S30)
);
Wallace w31(
	.n0(p0[31]),
	.n1(p1[31]),
	.n2(p2[31]),
	.n3(p3[31]),
	.n4(p4[31]),
	.n5(p5[31]),
	.n6(p6[31]),
	.n7(p7[31]),
	.n8(p8[31]),
	.n9(p9[31]),
	.n10(p10[31]),
	.n11(p11[31]),
	.n12(p12[31]),
	.n13(p13[31]),
	.n14(p14[31]),
	.n15(p15[31]),
	.cin0(cout30_0),
	.cin1(cout30_1),
	.cin2(cout30_2),
	.cin3(cout30_3),
	.cin4(cout30_4),
	.cin5(cout30_5),
	.cin6(cout30_6),
	.cin7(cout30_7),
	.cin8(cout30_8),
	.cin9(cout30_9),
	.cin10(cout30_10),
	.cin11(cout30_11),
	.cin12(cout30_12),
	.cin13(cout30_13),
	.c11(cout31_0),
	.c12(cout31_1),
	.c13(cout31_2),
	.c14(cout31_3),
	.c15(cout31_4),
	.c21(cout31_5),
	.c22(cout31_6),
	.c23(cout31_7),
	.c24(cout31_8),
	.c31(cout31_9),
	.c32(cout31_10),
	.c41(cout31_11),
	.c42(cout31_12),
	.c51(cout31_13),
	.c61(C31),
	.s61(S31)
);
Wallace w32(
	.n0(p0[32]),
	.n1(p1[32]),
	.n2(p2[32]),
	.n3(p3[32]),
	.n4(p4[32]),
	.n5(p5[32]),
	.n6(p6[32]),
	.n7(p7[32]),
	.n8(p8[32]),
	.n9(p9[32]),
	.n10(p10[32]),
	.n11(p11[32]),
	.n12(p12[32]),
	.n13(p13[32]),
	.n14(p14[32]),
	.n15(p15[32]),
	.cin0(cout31_0),
	.cin1(cout31_1),
	.cin2(cout31_2),
	.cin3(cout31_3),
	.cin4(cout31_4),
	.cin5(cout31_5),
	.cin6(cout31_6),
	.cin7(cout31_7),
	.cin8(cout31_8),
	.cin9(cout31_9),
	.cin10(cout31_10),
	.cin11(cout31_11),
	.cin12(cout31_12),
	.cin13(cout31_13),
	.c11(cout32_0),
	.c12(cout32_1),
	.c13(cout32_2),
	.c14(cout32_3),
	.c15(cout32_4),
	.c21(cout32_5),
	.c22(cout32_6),
	.c23(cout32_7),
	.c24(cout32_8),
	.c31(cout32_9),
	.c32(cout32_10),
	.c41(cout32_11),
	.c42(cout32_12),
	.c51(cout32_13),
	.c61(C32),
	.s61(S32)
);
Wallace w33(
	.n0(p0[33]),
	.n1(p1[33]),
	.n2(p2[33]),
	.n3(p3[33]),
	.n4(p4[33]),
	.n5(p5[33]),
	.n6(p6[33]),
	.n7(p7[33]),
	.n8(p8[33]),
	.n9(p9[33]),
	.n10(p10[33]),
	.n11(p11[33]),
	.n12(p12[33]),
	.n13(p13[33]),
	.n14(p14[33]),
	.n15(p15[33]),
	.cin0(cout32_0),
	.cin1(cout32_1),
	.cin2(cout32_2),
	.cin3(cout32_3),
	.cin4(cout32_4),
	.cin5(cout32_5),
	.cin6(cout32_6),
	.cin7(cout32_7),
	.cin8(cout32_8),
	.cin9(cout32_9),
	.cin10(cout32_10),
	.cin11(cout32_11),
	.cin12(cout32_12),
	.cin13(cout32_13),
	.c11(cout33_0),
	.c12(cout33_1),
	.c13(cout33_2),
	.c14(cout33_3),
	.c15(cout33_4),
	.c21(cout33_5),
	.c22(cout33_6),
	.c23(cout33_7),
	.c24(cout33_8),
	.c31(cout33_9),
	.c32(cout33_10),
	.c41(cout33_11),
	.c42(cout33_12),
	.c51(cout33_13),
	.c61(C33),
	.s61(S33)
);
Wallace w34(
	.n0(p0[34]),
	.n1(p1[34]),
	.n2(p2[34]),
	.n3(p3[34]),
	.n4(p4[34]),
	.n5(p5[34]),
	.n6(p6[34]),
	.n7(p7[34]),
	.n8(p8[34]),
	.n9(p9[34]),
	.n10(p10[34]),
	.n11(p11[34]),
	.n12(p12[34]),
	.n13(p13[34]),
	.n14(p14[34]),
	.n15(p15[34]),
	.cin0(cout33_0),
	.cin1(cout33_1),
	.cin2(cout33_2),
	.cin3(cout33_3),
	.cin4(cout33_4),
	.cin5(cout33_5),
	.cin6(cout33_6),
	.cin7(cout33_7),
	.cin8(cout33_8),
	.cin9(cout33_9),
	.cin10(cout33_10),
	.cin11(cout33_11),
	.cin12(cout33_12),
	.cin13(cout33_13),
	.c11(cout34_0),
	.c12(cout34_1),
	.c13(cout34_2),
	.c14(cout34_3),
	.c15(cout34_4),
	.c21(cout34_5),
	.c22(cout34_6),
	.c23(cout34_7),
	.c24(cout34_8),
	.c31(cout34_9),
	.c32(cout34_10),
	.c41(cout34_11),
	.c42(cout34_12),
	.c51(cout34_13),
	.c61(C34),
	.s61(S34)
);
Wallace w35(
	.n0(p0[35]),
	.n1(p1[35]),
	.n2(p2[35]),
	.n3(p3[35]),
	.n4(p4[35]),
	.n5(p5[35]),
	.n6(p6[35]),
	.n7(p7[35]),
	.n8(p8[35]),
	.n9(p9[35]),
	.n10(p10[35]),
	.n11(p11[35]),
	.n12(p12[35]),
	.n13(p13[35]),
	.n14(p14[35]),
	.n15(p15[35]),
	.cin0(cout34_0),
	.cin1(cout34_1),
	.cin2(cout34_2),
	.cin3(cout34_3),
	.cin4(cout34_4),
	.cin5(cout34_5),
	.cin6(cout34_6),
	.cin7(cout34_7),
	.cin8(cout34_8),
	.cin9(cout34_9),
	.cin10(cout34_10),
	.cin11(cout34_11),
	.cin12(cout34_12),
	.cin13(cout34_13),
	.c11(cout35_0),
	.c12(cout35_1),
	.c13(cout35_2),
	.c14(cout35_3),
	.c15(cout35_4),
	.c21(cout35_5),
	.c22(cout35_6),
	.c23(cout35_7),
	.c24(cout35_8),
	.c31(cout35_9),
	.c32(cout35_10),
	.c41(cout35_11),
	.c42(cout35_12),
	.c51(cout35_13),
	.c61(C35),
	.s61(S35)
);
Wallace w36(
	.n0(p0[36]),
	.n1(p1[36]),
	.n2(p2[36]),
	.n3(p3[36]),
	.n4(p4[36]),
	.n5(p5[36]),
	.n6(p6[36]),
	.n7(p7[36]),
	.n8(p8[36]),
	.n9(p9[36]),
	.n10(p10[36]),
	.n11(p11[36]),
	.n12(p12[36]),
	.n13(p13[36]),
	.n14(p14[36]),
	.n15(p15[36]),
	.cin0(cout35_0),
	.cin1(cout35_1),
	.cin2(cout35_2),
	.cin3(cout35_3),
	.cin4(cout35_4),
	.cin5(cout35_5),
	.cin6(cout35_6),
	.cin7(cout35_7),
	.cin8(cout35_8),
	.cin9(cout35_9),
	.cin10(cout35_10),
	.cin11(cout35_11),
	.cin12(cout35_12),
	.cin13(cout35_13),
	.c11(cout36_0),
	.c12(cout36_1),
	.c13(cout36_2),
	.c14(cout36_3),
	.c15(cout36_4),
	.c21(cout36_5),
	.c22(cout36_6),
	.c23(cout36_7),
	.c24(cout36_8),
	.c31(cout36_9),
	.c32(cout36_10),
	.c41(cout36_11),
	.c42(cout36_12),
	.c51(cout36_13),
	.c61(C36),
	.s61(S36)
);
Wallace w37(
	.n0(p0[37]),
	.n1(p1[37]),
	.n2(p2[37]),
	.n3(p3[37]),
	.n4(p4[37]),
	.n5(p5[37]),
	.n6(p6[37]),
	.n7(p7[37]),
	.n8(p8[37]),
	.n9(p9[37]),
	.n10(p10[37]),
	.n11(p11[37]),
	.n12(p12[37]),
	.n13(p13[37]),
	.n14(p14[37]),
	.n15(p15[37]),
	.cin0(cout36_0),
	.cin1(cout36_1),
	.cin2(cout36_2),
	.cin3(cout36_3),
	.cin4(cout36_4),
	.cin5(cout36_5),
	.cin6(cout36_6),
	.cin7(cout36_7),
	.cin8(cout36_8),
	.cin9(cout36_9),
	.cin10(cout36_10),
	.cin11(cout36_11),
	.cin12(cout36_12),
	.cin13(cout36_13),
	.c11(cout37_0),
	.c12(cout37_1),
	.c13(cout37_2),
	.c14(cout37_3),
	.c15(cout37_4),
	.c21(cout37_5),
	.c22(cout37_6),
	.c23(cout37_7),
	.c24(cout37_8),
	.c31(cout37_9),
	.c32(cout37_10),
	.c41(cout37_11),
	.c42(cout37_12),
	.c51(cout37_13),
	.c61(C37),
	.s61(S37)
);
Wallace w38(
	.n0(p0[38]),
	.n1(p1[38]),
	.n2(p2[38]),
	.n3(p3[38]),
	.n4(p4[38]),
	.n5(p5[38]),
	.n6(p6[38]),
	.n7(p7[38]),
	.n8(p8[38]),
	.n9(p9[38]),
	.n10(p10[38]),
	.n11(p11[38]),
	.n12(p12[38]),
	.n13(p13[38]),
	.n14(p14[38]),
	.n15(p15[38]),
	.cin0(cout37_0),
	.cin1(cout37_1),
	.cin2(cout37_2),
	.cin3(cout37_3),
	.cin4(cout37_4),
	.cin5(cout37_5),
	.cin6(cout37_6),
	.cin7(cout37_7),
	.cin8(cout37_8),
	.cin9(cout37_9),
	.cin10(cout37_10),
	.cin11(cout37_11),
	.cin12(cout37_12),
	.cin13(cout37_13),
	.c11(cout38_0),
	.c12(cout38_1),
	.c13(cout38_2),
	.c14(cout38_3),
	.c15(cout38_4),
	.c21(cout38_5),
	.c22(cout38_6),
	.c23(cout38_7),
	.c24(cout38_8),
	.c31(cout38_9),
	.c32(cout38_10),
	.c41(cout38_11),
	.c42(cout38_12),
	.c51(cout38_13),
	.c61(C38),
	.s61(S38)
);
Wallace w39(
	.n0(p0[39]),
	.n1(p1[39]),
	.n2(p2[39]),
	.n3(p3[39]),
	.n4(p4[39]),
	.n5(p5[39]),
	.n6(p6[39]),
	.n7(p7[39]),
	.n8(p8[39]),
	.n9(p9[39]),
	.n10(p10[39]),
	.n11(p11[39]),
	.n12(p12[39]),
	.n13(p13[39]),
	.n14(p14[39]),
	.n15(p15[39]),
	.cin0(cout38_0),
	.cin1(cout38_1),
	.cin2(cout38_2),
	.cin3(cout38_3),
	.cin4(cout38_4),
	.cin5(cout38_5),
	.cin6(cout38_6),
	.cin7(cout38_7),
	.cin8(cout38_8),
	.cin9(cout38_9),
	.cin10(cout38_10),
	.cin11(cout38_11),
	.cin12(cout38_12),
	.cin13(cout38_13),
	.c11(cout39_0),
	.c12(cout39_1),
	.c13(cout39_2),
	.c14(cout39_3),
	.c15(cout39_4),
	.c21(cout39_5),
	.c22(cout39_6),
	.c23(cout39_7),
	.c24(cout39_8),
	.c31(cout39_9),
	.c32(cout39_10),
	.c41(cout39_11),
	.c42(cout39_12),
	.c51(cout39_13),
	.c61(C39),
	.s61(S39)
);
Wallace w40(
	.n0(p0[40]),
	.n1(p1[40]),
	.n2(p2[40]),
	.n3(p3[40]),
	.n4(p4[40]),
	.n5(p5[40]),
	.n6(p6[40]),
	.n7(p7[40]),
	.n8(p8[40]),
	.n9(p9[40]),
	.n10(p10[40]),
	.n11(p11[40]),
	.n12(p12[40]),
	.n13(p13[40]),
	.n14(p14[40]),
	.n15(p15[40]),
	.cin0(cout39_0),
	.cin1(cout39_1),
	.cin2(cout39_2),
	.cin3(cout39_3),
	.cin4(cout39_4),
	.cin5(cout39_5),
	.cin6(cout39_6),
	.cin7(cout39_7),
	.cin8(cout39_8),
	.cin9(cout39_9),
	.cin10(cout39_10),
	.cin11(cout39_11),
	.cin12(cout39_12),
	.cin13(cout39_13),
	.c11(cout40_0),
	.c12(cout40_1),
	.c13(cout40_2),
	.c14(cout40_3),
	.c15(cout40_4),
	.c21(cout40_5),
	.c22(cout40_6),
	.c23(cout40_7),
	.c24(cout40_8),
	.c31(cout40_9),
	.c32(cout40_10),
	.c41(cout40_11),
	.c42(cout40_12),
	.c51(cout40_13),
	.c61(C40),
	.s61(S40)
);
Wallace w41(
	.n0(p0[41]),
	.n1(p1[41]),
	.n2(p2[41]),
	.n3(p3[41]),
	.n4(p4[41]),
	.n5(p5[41]),
	.n6(p6[41]),
	.n7(p7[41]),
	.n8(p8[41]),
	.n9(p9[41]),
	.n10(p10[41]),
	.n11(p11[41]),
	.n12(p12[41]),
	.n13(p13[41]),
	.n14(p14[41]),
	.n15(p15[41]),
	.cin0(cout40_0),
	.cin1(cout40_1),
	.cin2(cout40_2),
	.cin3(cout40_3),
	.cin4(cout40_4),
	.cin5(cout40_5),
	.cin6(cout40_6),
	.cin7(cout40_7),
	.cin8(cout40_8),
	.cin9(cout40_9),
	.cin10(cout40_10),
	.cin11(cout40_11),
	.cin12(cout40_12),
	.cin13(cout40_13),
	.c11(cout41_0),
	.c12(cout41_1),
	.c13(cout41_2),
	.c14(cout41_3),
	.c15(cout41_4),
	.c21(cout41_5),
	.c22(cout41_6),
	.c23(cout41_7),
	.c24(cout41_8),
	.c31(cout41_9),
	.c32(cout41_10),
	.c41(cout41_11),
	.c42(cout41_12),
	.c51(cout41_13),
	.c61(C41),
	.s61(S41)
);
Wallace w42(
	.n0(p0[42]),
	.n1(p1[42]),
	.n2(p2[42]),
	.n3(p3[42]),
	.n4(p4[42]),
	.n5(p5[42]),
	.n6(p6[42]),
	.n7(p7[42]),
	.n8(p8[42]),
	.n9(p9[42]),
	.n10(p10[42]),
	.n11(p11[42]),
	.n12(p12[42]),
	.n13(p13[42]),
	.n14(p14[42]),
	.n15(p15[42]),
	.cin0(cout41_0),
	.cin1(cout41_1),
	.cin2(cout41_2),
	.cin3(cout41_3),
	.cin4(cout41_4),
	.cin5(cout41_5),
	.cin6(cout41_6),
	.cin7(cout41_7),
	.cin8(cout41_8),
	.cin9(cout41_9),
	.cin10(cout41_10),
	.cin11(cout41_11),
	.cin12(cout41_12),
	.cin13(cout41_13),
	.c11(cout42_0),
	.c12(cout42_1),
	.c13(cout42_2),
	.c14(cout42_3),
	.c15(cout42_4),
	.c21(cout42_5),
	.c22(cout42_6),
	.c23(cout42_7),
	.c24(cout42_8),
	.c31(cout42_9),
	.c32(cout42_10),
	.c41(cout42_11),
	.c42(cout42_12),
	.c51(cout42_13),
	.c61(C42),
	.s61(S42)
);
Wallace w43(
	.n0(p0[43]),
	.n1(p1[43]),
	.n2(p2[43]),
	.n3(p3[43]),
	.n4(p4[43]),
	.n5(p5[43]),
	.n6(p6[43]),
	.n7(p7[43]),
	.n8(p8[43]),
	.n9(p9[43]),
	.n10(p10[43]),
	.n11(p11[43]),
	.n12(p12[43]),
	.n13(p13[43]),
	.n14(p14[43]),
	.n15(p15[43]),
	.cin0(cout42_0),
	.cin1(cout42_1),
	.cin2(cout42_2),
	.cin3(cout42_3),
	.cin4(cout42_4),
	.cin5(cout42_5),
	.cin6(cout42_6),
	.cin7(cout42_7),
	.cin8(cout42_8),
	.cin9(cout42_9),
	.cin10(cout42_10),
	.cin11(cout42_11),
	.cin12(cout42_12),
	.cin13(cout42_13),
	.c11(cout43_0),
	.c12(cout43_1),
	.c13(cout43_2),
	.c14(cout43_3),
	.c15(cout43_4),
	.c21(cout43_5),
	.c22(cout43_6),
	.c23(cout43_7),
	.c24(cout43_8),
	.c31(cout43_9),
	.c32(cout43_10),
	.c41(cout43_11),
	.c42(cout43_12),
	.c51(cout43_13),
	.c61(C43),
	.s61(S43)
);
Wallace w44(
	.n0(p0[44]),
	.n1(p1[44]),
	.n2(p2[44]),
	.n3(p3[44]),
	.n4(p4[44]),
	.n5(p5[44]),
	.n6(p6[44]),
	.n7(p7[44]),
	.n8(p8[44]),
	.n9(p9[44]),
	.n10(p10[44]),
	.n11(p11[44]),
	.n12(p12[44]),
	.n13(p13[44]),
	.n14(p14[44]),
	.n15(p15[44]),
	.cin0(cout43_0),
	.cin1(cout43_1),
	.cin2(cout43_2),
	.cin3(cout43_3),
	.cin4(cout43_4),
	.cin5(cout43_5),
	.cin6(cout43_6),
	.cin7(cout43_7),
	.cin8(cout43_8),
	.cin9(cout43_9),
	.cin10(cout43_10),
	.cin11(cout43_11),
	.cin12(cout43_12),
	.cin13(cout43_13),
	.c11(cout44_0),
	.c12(cout44_1),
	.c13(cout44_2),
	.c14(cout44_3),
	.c15(cout44_4),
	.c21(cout44_5),
	.c22(cout44_6),
	.c23(cout44_7),
	.c24(cout44_8),
	.c31(cout44_9),
	.c32(cout44_10),
	.c41(cout44_11),
	.c42(cout44_12),
	.c51(cout44_13),
	.c61(C44),
	.s61(S44)
);
Wallace w45(
	.n0(p0[45]),
	.n1(p1[45]),
	.n2(p2[45]),
	.n3(p3[45]),
	.n4(p4[45]),
	.n5(p5[45]),
	.n6(p6[45]),
	.n7(p7[45]),
	.n8(p8[45]),
	.n9(p9[45]),
	.n10(p10[45]),
	.n11(p11[45]),
	.n12(p12[45]),
	.n13(p13[45]),
	.n14(p14[45]),
	.n15(p15[45]),
	.cin0(cout44_0),
	.cin1(cout44_1),
	.cin2(cout44_2),
	.cin3(cout44_3),
	.cin4(cout44_4),
	.cin5(cout44_5),
	.cin6(cout44_6),
	.cin7(cout44_7),
	.cin8(cout44_8),
	.cin9(cout44_9),
	.cin10(cout44_10),
	.cin11(cout44_11),
	.cin12(cout44_12),
	.cin13(cout44_13),
	.c11(cout45_0),
	.c12(cout45_1),
	.c13(cout45_2),
	.c14(cout45_3),
	.c15(cout45_4),
	.c21(cout45_5),
	.c22(cout45_6),
	.c23(cout45_7),
	.c24(cout45_8),
	.c31(cout45_9),
	.c32(cout45_10),
	.c41(cout45_11),
	.c42(cout45_12),
	.c51(cout45_13),
	.c61(C45),
	.s61(S45)
);
Wallace w46(
	.n0(p0[46]),
	.n1(p1[46]),
	.n2(p2[46]),
	.n3(p3[46]),
	.n4(p4[46]),
	.n5(p5[46]),
	.n6(p6[46]),
	.n7(p7[46]),
	.n8(p8[46]),
	.n9(p9[46]),
	.n10(p10[46]),
	.n11(p11[46]),
	.n12(p12[46]),
	.n13(p13[46]),
	.n14(p14[46]),
	.n15(p15[46]),
	.cin0(cout45_0),
	.cin1(cout45_1),
	.cin2(cout45_2),
	.cin3(cout45_3),
	.cin4(cout45_4),
	.cin5(cout45_5),
	.cin6(cout45_6),
	.cin7(cout45_7),
	.cin8(cout45_8),
	.cin9(cout45_9),
	.cin10(cout45_10),
	.cin11(cout45_11),
	.cin12(cout45_12),
	.cin13(cout45_13),
	.c11(cout46_0),
	.c12(cout46_1),
	.c13(cout46_2),
	.c14(cout46_3),
	.c15(cout46_4),
	.c21(cout46_5),
	.c22(cout46_6),
	.c23(cout46_7),
	.c24(cout46_8),
	.c31(cout46_9),
	.c32(cout46_10),
	.c41(cout46_11),
	.c42(cout46_12),
	.c51(cout46_13),
	.c61(C46),
	.s61(S46)
);
Wallace w47(
	.n0(p0[47]),
	.n1(p1[47]),
	.n2(p2[47]),
	.n3(p3[47]),
	.n4(p4[47]),
	.n5(p5[47]),
	.n6(p6[47]),
	.n7(p7[47]),
	.n8(p8[47]),
	.n9(p9[47]),
	.n10(p10[47]),
	.n11(p11[47]),
	.n12(p12[47]),
	.n13(p13[47]),
	.n14(p14[47]),
	.n15(p15[47]),
	.cin0(cout46_0),
	.cin1(cout46_1),
	.cin2(cout46_2),
	.cin3(cout46_3),
	.cin4(cout46_4),
	.cin5(cout46_5),
	.cin6(cout46_6),
	.cin7(cout46_7),
	.cin8(cout46_8),
	.cin9(cout46_9),
	.cin10(cout46_10),
	.cin11(cout46_11),
	.cin12(cout46_12),
	.cin13(cout46_13),
	.c11(cout47_0),
	.c12(cout47_1),
	.c13(cout47_2),
	.c14(cout47_3),
	.c15(cout47_4),
	.c21(cout47_5),
	.c22(cout47_6),
	.c23(cout47_7),
	.c24(cout47_8),
	.c31(cout47_9),
	.c32(cout47_10),
	.c41(cout47_11),
	.c42(cout47_12),
	.c51(cout47_13),
	.c61(C47),
	.s61(S47)
);
Wallace w48(
	.n0(p0[48]),
	.n1(p1[48]),
	.n2(p2[48]),
	.n3(p3[48]),
	.n4(p4[48]),
	.n5(p5[48]),
	.n6(p6[48]),
	.n7(p7[48]),
	.n8(p8[48]),
	.n9(p9[48]),
	.n10(p10[48]),
	.n11(p11[48]),
	.n12(p12[48]),
	.n13(p13[48]),
	.n14(p14[48]),
	.n15(p15[48]),
	.cin0(cout47_0),
	.cin1(cout47_1),
	.cin2(cout47_2),
	.cin3(cout47_3),
	.cin4(cout47_4),
	.cin5(cout47_5),
	.cin6(cout47_6),
	.cin7(cout47_7),
	.cin8(cout47_8),
	.cin9(cout47_9),
	.cin10(cout47_10),
	.cin11(cout47_11),
	.cin12(cout47_12),
	.cin13(cout47_13),
	.c11(cout48_0),
	.c12(cout48_1),
	.c13(cout48_2),
	.c14(cout48_3),
	.c15(cout48_4),
	.c21(cout48_5),
	.c22(cout48_6),
	.c23(cout48_7),
	.c24(cout48_8),
	.c31(cout48_9),
	.c32(cout48_10),
	.c41(cout48_11),
	.c42(cout48_12),
	.c51(cout48_13),
	.c61(C48),
	.s61(S48)
);
Wallace w49(
	.n0(p0[49]),
	.n1(p1[49]),
	.n2(p2[49]),
	.n3(p3[49]),
	.n4(p4[49]),
	.n5(p5[49]),
	.n6(p6[49]),
	.n7(p7[49]),
	.n8(p8[49]),
	.n9(p9[49]),
	.n10(p10[49]),
	.n11(p11[49]),
	.n12(p12[49]),
	.n13(p13[49]),
	.n14(p14[49]),
	.n15(p15[49]),
	.cin0(cout48_0),
	.cin1(cout48_1),
	.cin2(cout48_2),
	.cin3(cout48_3),
	.cin4(cout48_4),
	.cin5(cout48_5),
	.cin6(cout48_6),
	.cin7(cout48_7),
	.cin8(cout48_8),
	.cin9(cout48_9),
	.cin10(cout48_10),
	.cin11(cout48_11),
	.cin12(cout48_12),
	.cin13(cout48_13),
	.c11(cout49_0),
	.c12(cout49_1),
	.c13(cout49_2),
	.c14(cout49_3),
	.c15(cout49_4),
	.c21(cout49_5),
	.c22(cout49_6),
	.c23(cout49_7),
	.c24(cout49_8),
	.c31(cout49_9),
	.c32(cout49_10),
	.c41(cout49_11),
	.c42(cout49_12),
	.c51(cout49_13),
	.c61(C49),
	.s61(S49)
);
Wallace w50(
	.n0(p0[50]),
	.n1(p1[50]),
	.n2(p2[50]),
	.n3(p3[50]),
	.n4(p4[50]),
	.n5(p5[50]),
	.n6(p6[50]),
	.n7(p7[50]),
	.n8(p8[50]),
	.n9(p9[50]),
	.n10(p10[50]),
	.n11(p11[50]),
	.n12(p12[50]),
	.n13(p13[50]),
	.n14(p14[50]),
	.n15(p15[50]),
	.cin0(cout49_0),
	.cin1(cout49_1),
	.cin2(cout49_2),
	.cin3(cout49_3),
	.cin4(cout49_4),
	.cin5(cout49_5),
	.cin6(cout49_6),
	.cin7(cout49_7),
	.cin8(cout49_8),
	.cin9(cout49_9),
	.cin10(cout49_10),
	.cin11(cout49_11),
	.cin12(cout49_12),
	.cin13(cout49_13),
	.c11(cout50_0),
	.c12(cout50_1),
	.c13(cout50_2),
	.c14(cout50_3),
	.c15(cout50_4),
	.c21(cout50_5),
	.c22(cout50_6),
	.c23(cout50_7),
	.c24(cout50_8),
	.c31(cout50_9),
	.c32(cout50_10),
	.c41(cout50_11),
	.c42(cout50_12),
	.c51(cout50_13),
	.c61(C50),
	.s61(S50)
);
Wallace w51(
	.n0(p0[51]),
	.n1(p1[51]),
	.n2(p2[51]),
	.n3(p3[51]),
	.n4(p4[51]),
	.n5(p5[51]),
	.n6(p6[51]),
	.n7(p7[51]),
	.n8(p8[51]),
	.n9(p9[51]),
	.n10(p10[51]),
	.n11(p11[51]),
	.n12(p12[51]),
	.n13(p13[51]),
	.n14(p14[51]),
	.n15(p15[51]),
	.cin0(cout50_0),
	.cin1(cout50_1),
	.cin2(cout50_2),
	.cin3(cout50_3),
	.cin4(cout50_4),
	.cin5(cout50_5),
	.cin6(cout50_6),
	.cin7(cout50_7),
	.cin8(cout50_8),
	.cin9(cout50_9),
	.cin10(cout50_10),
	.cin11(cout50_11),
	.cin12(cout50_12),
	.cin13(cout50_13),
	.c11(cout51_0),
	.c12(cout51_1),
	.c13(cout51_2),
	.c14(cout51_3),
	.c15(cout51_4),
	.c21(cout51_5),
	.c22(cout51_6),
	.c23(cout51_7),
	.c24(cout51_8),
	.c31(cout51_9),
	.c32(cout51_10),
	.c41(cout51_11),
	.c42(cout51_12),
	.c51(cout51_13),
	.c61(C51),
	.s61(S51)
);
Wallace w52(
	.n0(p0[52]),
	.n1(p1[52]),
	.n2(p2[52]),
	.n3(p3[52]),
	.n4(p4[52]),
	.n5(p5[52]),
	.n6(p6[52]),
	.n7(p7[52]),
	.n8(p8[52]),
	.n9(p9[52]),
	.n10(p10[52]),
	.n11(p11[52]),
	.n12(p12[52]),
	.n13(p13[52]),
	.n14(p14[52]),
	.n15(p15[52]),
	.cin0(cout51_0),
	.cin1(cout51_1),
	.cin2(cout51_2),
	.cin3(cout51_3),
	.cin4(cout51_4),
	.cin5(cout51_5),
	.cin6(cout51_6),
	.cin7(cout51_7),
	.cin8(cout51_8),
	.cin9(cout51_9),
	.cin10(cout51_10),
	.cin11(cout51_11),
	.cin12(cout51_12),
	.cin13(cout51_13),
	.c11(cout52_0),
	.c12(cout52_1),
	.c13(cout52_2),
	.c14(cout52_3),
	.c15(cout52_4),
	.c21(cout52_5),
	.c22(cout52_6),
	.c23(cout52_7),
	.c24(cout52_8),
	.c31(cout52_9),
	.c32(cout52_10),
	.c41(cout52_11),
	.c42(cout52_12),
	.c51(cout52_13),
	.c61(C52),
	.s61(S52)
);
Wallace w53(
	.n0(p0[53]),
	.n1(p1[53]),
	.n2(p2[53]),
	.n3(p3[53]),
	.n4(p4[53]),
	.n5(p5[53]),
	.n6(p6[53]),
	.n7(p7[53]),
	.n8(p8[53]),
	.n9(p9[53]),
	.n10(p10[53]),
	.n11(p11[53]),
	.n12(p12[53]),
	.n13(p13[53]),
	.n14(p14[53]),
	.n15(p15[53]),
	.cin0(cout52_0),
	.cin1(cout52_1),
	.cin2(cout52_2),
	.cin3(cout52_3),
	.cin4(cout52_4),
	.cin5(cout52_5),
	.cin6(cout52_6),
	.cin7(cout52_7),
	.cin8(cout52_8),
	.cin9(cout52_9),
	.cin10(cout52_10),
	.cin11(cout52_11),
	.cin12(cout52_12),
	.cin13(cout52_13),
	.c11(cout53_0),
	.c12(cout53_1),
	.c13(cout53_2),
	.c14(cout53_3),
	.c15(cout53_4),
	.c21(cout53_5),
	.c22(cout53_6),
	.c23(cout53_7),
	.c24(cout53_8),
	.c31(cout53_9),
	.c32(cout53_10),
	.c41(cout53_11),
	.c42(cout53_12),
	.c51(cout53_13),
	.c61(C53),
	.s61(S53)
);
Wallace w54(
	.n0(p0[54]),
	.n1(p1[54]),
	.n2(p2[54]),
	.n3(p3[54]),
	.n4(p4[54]),
	.n5(p5[54]),
	.n6(p6[54]),
	.n7(p7[54]),
	.n8(p8[54]),
	.n9(p9[54]),
	.n10(p10[54]),
	.n11(p11[54]),
	.n12(p12[54]),
	.n13(p13[54]),
	.n14(p14[54]),
	.n15(p15[54]),
	.cin0(cout53_0),
	.cin1(cout53_1),
	.cin2(cout53_2),
	.cin3(cout53_3),
	.cin4(cout53_4),
	.cin5(cout53_5),
	.cin6(cout53_6),
	.cin7(cout53_7),
	.cin8(cout53_8),
	.cin9(cout53_9),
	.cin10(cout53_10),
	.cin11(cout53_11),
	.cin12(cout53_12),
	.cin13(cout53_13),
	.c11(cout54_0),
	.c12(cout54_1),
	.c13(cout54_2),
	.c14(cout54_3),
	.c15(cout54_4),
	.c21(cout54_5),
	.c22(cout54_6),
	.c23(cout54_7),
	.c24(cout54_8),
	.c31(cout54_9),
	.c32(cout54_10),
	.c41(cout54_11),
	.c42(cout54_12),
	.c51(cout54_13),
	.c61(C54),
	.s61(S54)
);
Wallace w55(
	.n0(p0[55]),
	.n1(p1[55]),
	.n2(p2[55]),
	.n3(p3[55]),
	.n4(p4[55]),
	.n5(p5[55]),
	.n6(p6[55]),
	.n7(p7[55]),
	.n8(p8[55]),
	.n9(p9[55]),
	.n10(p10[55]),
	.n11(p11[55]),
	.n12(p12[55]),
	.n13(p13[55]),
	.n14(p14[55]),
	.n15(p15[55]),
	.cin0(cout54_0),
	.cin1(cout54_1),
	.cin2(cout54_2),
	.cin3(cout54_3),
	.cin4(cout54_4),
	.cin5(cout54_5),
	.cin6(cout54_6),
	.cin7(cout54_7),
	.cin8(cout54_8),
	.cin9(cout54_9),
	.cin10(cout54_10),
	.cin11(cout54_11),
	.cin12(cout54_12),
	.cin13(cout54_13),
	.c11(cout55_0),
	.c12(cout55_1),
	.c13(cout55_2),
	.c14(cout55_3),
	.c15(cout55_4),
	.c21(cout55_5),
	.c22(cout55_6),
	.c23(cout55_7),
	.c24(cout55_8),
	.c31(cout55_9),
	.c32(cout55_10),
	.c41(cout55_11),
	.c42(cout55_12),
	.c51(cout55_13),
	.c61(C55),
	.s61(S55)
);
Wallace w56(
	.n0(p0[56]),
	.n1(p1[56]),
	.n2(p2[56]),
	.n3(p3[56]),
	.n4(p4[56]),
	.n5(p5[56]),
	.n6(p6[56]),
	.n7(p7[56]),
	.n8(p8[56]),
	.n9(p9[56]),
	.n10(p10[56]),
	.n11(p11[56]),
	.n12(p12[56]),
	.n13(p13[56]),
	.n14(p14[56]),
	.n15(p15[56]),
	.cin0(cout55_0),
	.cin1(cout55_1),
	.cin2(cout55_2),
	.cin3(cout55_3),
	.cin4(cout55_4),
	.cin5(cout55_5),
	.cin6(cout55_6),
	.cin7(cout55_7),
	.cin8(cout55_8),
	.cin9(cout55_9),
	.cin10(cout55_10),
	.cin11(cout55_11),
	.cin12(cout55_12),
	.cin13(cout55_13),
	.c11(cout56_0),
	.c12(cout56_1),
	.c13(cout56_2),
	.c14(cout56_3),
	.c15(cout56_4),
	.c21(cout56_5),
	.c22(cout56_6),
	.c23(cout56_7),
	.c24(cout56_8),
	.c31(cout56_9),
	.c32(cout56_10),
	.c41(cout56_11),
	.c42(cout56_12),
	.c51(cout56_13),
	.c61(C56),
	.s61(S56)
);
Wallace w57(
	.n0(p0[57]),
	.n1(p1[57]),
	.n2(p2[57]),
	.n3(p3[57]),
	.n4(p4[57]),
	.n5(p5[57]),
	.n6(p6[57]),
	.n7(p7[57]),
	.n8(p8[57]),
	.n9(p9[57]),
	.n10(p10[57]),
	.n11(p11[57]),
	.n12(p12[57]),
	.n13(p13[57]),
	.n14(p14[57]),
	.n15(p15[57]),
	.cin0(cout56_0),
	.cin1(cout56_1),
	.cin2(cout56_2),
	.cin3(cout56_3),
	.cin4(cout56_4),
	.cin5(cout56_5),
	.cin6(cout56_6),
	.cin7(cout56_7),
	.cin8(cout56_8),
	.cin9(cout56_9),
	.cin10(cout56_10),
	.cin11(cout56_11),
	.cin12(cout56_12),
	.cin13(cout56_13),
	.c11(cout57_0),
	.c12(cout57_1),
	.c13(cout57_2),
	.c14(cout57_3),
	.c15(cout57_4),
	.c21(cout57_5),
	.c22(cout57_6),
	.c23(cout57_7),
	.c24(cout57_8),
	.c31(cout57_9),
	.c32(cout57_10),
	.c41(cout57_11),
	.c42(cout57_12),
	.c51(cout57_13),
	.c61(C57),
	.s61(S57)
);
Wallace w58(
	.n0(p0[58]),
	.n1(p1[58]),
	.n2(p2[58]),
	.n3(p3[58]),
	.n4(p4[58]),
	.n5(p5[58]),
	.n6(p6[58]),
	.n7(p7[58]),
	.n8(p8[58]),
	.n9(p9[58]),
	.n10(p10[58]),
	.n11(p11[58]),
	.n12(p12[58]),
	.n13(p13[58]),
	.n14(p14[58]),
	.n15(p15[58]),
	.cin0(cout57_0),
	.cin1(cout57_1),
	.cin2(cout57_2),
	.cin3(cout57_3),
	.cin4(cout57_4),
	.cin5(cout57_5),
	.cin6(cout57_6),
	.cin7(cout57_7),
	.cin8(cout57_8),
	.cin9(cout57_9),
	.cin10(cout57_10),
	.cin11(cout57_11),
	.cin12(cout57_12),
	.cin13(cout57_13),
	.c11(cout58_0),
	.c12(cout58_1),
	.c13(cout58_2),
	.c14(cout58_3),
	.c15(cout58_4),
	.c21(cout58_5),
	.c22(cout58_6),
	.c23(cout58_7),
	.c24(cout58_8),
	.c31(cout58_9),
	.c32(cout58_10),
	.c41(cout58_11),
	.c42(cout58_12),
	.c51(cout58_13),
	.c61(C58),
	.s61(S58)
);
Wallace w59(
	.n0(p0[59]),
	.n1(p1[59]),
	.n2(p2[59]),
	.n3(p3[59]),
	.n4(p4[59]),
	.n5(p5[59]),
	.n6(p6[59]),
	.n7(p7[59]),
	.n8(p8[59]),
	.n9(p9[59]),
	.n10(p10[59]),
	.n11(p11[59]),
	.n12(p12[59]),
	.n13(p13[59]),
	.n14(p14[59]),
	.n15(p15[59]),
	.cin0(cout58_0),
	.cin1(cout58_1),
	.cin2(cout58_2),
	.cin3(cout58_3),
	.cin4(cout58_4),
	.cin5(cout58_5),
	.cin6(cout58_6),
	.cin7(cout58_7),
	.cin8(cout58_8),
	.cin9(cout58_9),
	.cin10(cout58_10),
	.cin11(cout58_11),
	.cin12(cout58_12),
	.cin13(cout58_13),
	.c11(cout59_0),
	.c12(cout59_1),
	.c13(cout59_2),
	.c14(cout59_3),
	.c15(cout59_4),
	.c21(cout59_5),
	.c22(cout59_6),
	.c23(cout59_7),
	.c24(cout59_8),
	.c31(cout59_9),
	.c32(cout59_10),
	.c41(cout59_11),
	.c42(cout59_12),
	.c51(cout59_13),
	.c61(C59),
	.s61(S59)
);
Wallace w60(
	.n0(p0[60]),
	.n1(p1[60]),
	.n2(p2[60]),
	.n3(p3[60]),
	.n4(p4[60]),
	.n5(p5[60]),
	.n6(p6[60]),
	.n7(p7[60]),
	.n8(p8[60]),
	.n9(p9[60]),
	.n10(p10[60]),
	.n11(p11[60]),
	.n12(p12[60]),
	.n13(p13[60]),
	.n14(p14[60]),
	.n15(p15[60]),
	.cin0(cout59_0),
	.cin1(cout59_1),
	.cin2(cout59_2),
	.cin3(cout59_3),
	.cin4(cout59_4),
	.cin5(cout59_5),
	.cin6(cout59_6),
	.cin7(cout59_7),
	.cin8(cout59_8),
	.cin9(cout59_9),
	.cin10(cout59_10),
	.cin11(cout59_11),
	.cin12(cout59_12),
	.cin13(cout59_13),
	.c11(cout60_0),
	.c12(cout60_1),
	.c13(cout60_2),
	.c14(cout60_3),
	.c15(cout60_4),
	.c21(cout60_5),
	.c22(cout60_6),
	.c23(cout60_7),
	.c24(cout60_8),
	.c31(cout60_9),
	.c32(cout60_10),
	.c41(cout60_11),
	.c42(cout60_12),
	.c51(cout60_13),
	.c61(C60),
	.s61(S60)
);
Wallace w61(
	.n0(p0[61]),
	.n1(p1[61]),
	.n2(p2[61]),
	.n3(p3[61]),
	.n4(p4[61]),
	.n5(p5[61]),
	.n6(p6[61]),
	.n7(p7[61]),
	.n8(p8[61]),
	.n9(p9[61]),
	.n10(p10[61]),
	.n11(p11[61]),
	.n12(p12[61]),
	.n13(p13[61]),
	.n14(p14[61]),
	.n15(p15[61]),
	.cin0(cout60_0),
	.cin1(cout60_1),
	.cin2(cout60_2),
	.cin3(cout60_3),
	.cin4(cout60_4),
	.cin5(cout60_5),
	.cin6(cout60_6),
	.cin7(cout60_7),
	.cin8(cout60_8),
	.cin9(cout60_9),
	.cin10(cout60_10),
	.cin11(cout60_11),
	.cin12(cout60_12),
	.cin13(cout60_13),
	.c11(cout61_0),
	.c12(cout61_1),
	.c13(cout61_2),
	.c14(cout61_3),
	.c15(cout61_4),
	.c21(cout61_5),
	.c22(cout61_6),
	.c23(cout61_7),
	.c24(cout61_8),
	.c31(cout61_9),
	.c32(cout61_10),
	.c41(cout61_11),
	.c42(cout61_12),
	.c51(cout61_13),
	.c61(C61),
	.s61(S61)
);
Wallace w62(
	.n0(p0[62]),
	.n1(p1[62]),
	.n2(p2[62]),
	.n3(p3[62]),
	.n4(p4[62]),
	.n5(p5[62]),
	.n6(p6[62]),
	.n7(p7[62]),
	.n8(p8[62]),
	.n9(p9[62]),
	.n10(p10[62]),
	.n11(p11[62]),
	.n12(p12[62]),
	.n13(p13[62]),
	.n14(p14[62]),
	.n15(p15[62]),
	.cin0(cout61_0),
	.cin1(cout61_1),
	.cin2(cout61_2),
	.cin3(cout61_3),
	.cin4(cout61_4),
	.cin5(cout61_5),
	.cin6(cout61_6),
	.cin7(cout61_7),
	.cin8(cout61_8),
	.cin9(cout61_9),
	.cin10(cout61_10),
	.cin11(cout61_11),
	.cin12(cout61_12),
	.cin13(cout61_13),
	.c11(cout62_0),
	.c12(cout62_1),
	.c13(cout62_2),
	.c14(cout62_3),
	.c15(cout62_4),
	.c21(cout62_5),
	.c22(cout62_6),
	.c23(cout62_7),
	.c24(cout62_8),
	.c31(cout62_9),
	.c32(cout62_10),
	.c41(cout62_11),
	.c42(cout62_12),
	.c51(cout62_13),
	.c61(C62),
	.s61(S62)
);
Wallace w63(
	.n0(p0[63]),
	.n1(p1[63]),
	.n2(p2[63]),
	.n3(p3[63]),
	.n4(p4[63]),
	.n5(p5[63]),
	.n6(p6[63]),
	.n7(p7[63]),
	.n8(p8[63]),
	.n9(p9[63]),
	.n10(p10[63]),
	.n11(p11[63]),
	.n12(p12[63]),
	.n13(p13[63]),
	.n14(p14[63]),
	.n15(p15[63]),
	.cin0(cout62_0),
	.cin1(cout62_1),
	.cin2(cout62_2),
	.cin3(cout62_3),
	.cin4(cout62_4),
	.cin5(cout62_5),
	.cin6(cout62_6),
	.cin7(cout62_7),
	.cin8(cout62_8),
	.cin9(cout62_9),
	.cin10(cout62_10),
	.cin11(cout62_11),
	.cin12(cout62_12),
	.cin13(cout62_13),
	.c11(cout63_0),
	.c12(cout63_1),
	.c13(cout63_2),
	.c14(cout63_3),
	.c15(cout63_4),
	.c21(cout63_5),
	.c22(cout63_6),
	.c23(cout63_7),
	.c24(cout63_8),
	.c31(cout63_9),
	.c32(cout63_10),
	.c41(cout63_11),
	.c42(cout63_12),
	.c51(cout63_13),
	.c61(C63),
	.s61(S63)
);

endmodule

module booth(
    input y2,
    input y1,
    input y0,
    input [63:0] X,
    output [63:0] p,
    output c
);

wire addx,add2x,subx,sub2x;
assign addx = ~y2&y1&~y0|~y2&~y1&y0;
assign add2x = ~y2&y1&y0;
assign subx = y2&y1&~y0|y2&~y1&y0;
assign sub2x = y2&~y1&~y0;
assign c = subx | sub2x;
assign p[0] = subx&~X[0] | addx&X[0] | sub2x;
genvar nbit;
generate 
    for(nbit = 1; nbit<64; nbit = nbit+1)
        begin: kkk
            assign p[nbit] = subx&~X[nbit]|sub2x&~X[nbit-1]|addx&X[nbit]|add2x&X[nbit-1];
        end
    
endgenerate

endmodule

module Full_adder(
    input A,
    input B,
    input cin,
    output sum,
    output cout
);
assign sum = ~A & ~B & cin | ~A & B & ~cin | A & ~B & ~cin | A & B & cin;
assign cout = A & B | A & cin | B & cin;

endmodule

module Wallace(
    input n0,
    input n1,
    input n2,
    input n3,
    input n4,
    input n5,
    input n6,
    input n7,
    input n8,
    input n9,
    input n10,
    input n11,
    input n12,
    input n13,
    input n14,
    input n15,
    input cin0,
    input cin1,
    input cin2,
    input cin3,
    input cin4,
    input cin5,
    input cin6,
    input cin7,
    input cin8,
    input cin9,
    input cin10,
    input cin11,
    input cin12,
    input cin13,
    output c11,
    output c12,
    output c13,
    output c14,
    output c15,
    output c21,
    output c22,
    output c23,
    output c24,
    output c31,
    output c32,
    output c41,
    output c42,
    output c51,
    output c61,
    output s61
);
wire s11,s12,s13,s14,s15;
wire s21,s22,s23,s24;
wire s31,s32;
wire s41,s42;
wire s51;

Full_adder a11(
    .A(n0),
    .B(n1),
    .cin(n2),
    .sum(s11),
    .cout(c11)
);
Full_adder a12(
    .A(n3),
    .B(n4),
    .cin(n5),
    .sum(s12),
    .cout(c12)
);
Full_adder a13(
    .A(n6),
    .B(n7),
    .cin(n8),
    .sum(s13),
    .cout(c13)
);
Full_adder a14(
    .A(n9),
    .B(n10),
    .cin(n11),
    .sum(s14),
    .cout(c14)
);
Full_adder a15(
    .A(n12),
    .B(n13),
    .cin(n14),
    .sum(s15),
    .cout(c15)
);
Full_adder a21(
    .A(s11),
    .B(s12),
    .cin(s13),
    .sum(s21),
    .cout(c21)
);
Full_adder a22(
    .A(s14),
    .B(s15),
    .cin(n15),
    .sum(s22),
    .cout(c22)
);
Full_adder a23(
    .A(cin0),
    .B(cin1),
    .cin(cin2),
    .sum(s23),
    .cout(c23)
);
Full_adder a24(
    .A(cin3),
    .B(cin4),
    .cin(0),
    .sum(s24),
    .cout(c24)
);
Full_adder a31(
    .A(s21),
    .B(s22),
    .cin(s23),
    .sum(s31),
    .cout(c31)
);
Full_adder a32(
    .A(s24),
    .B(cin5),
    .cin(cin6),
    .sum(s32),
    .cout(c32)
);
Full_adder a41(
    .A(s31),
    .B(s32),
    .cin(cin7),
    .sum(s41),
    .cout(c41)
);
Full_adder a42(
    .A(cin8),
    .B(cin9),
    .cin(cin10),
    .sum(s42),
    .cout(c42)
);
Full_adder a51(
    .A(s41),
    .B(s42),
    .cin(cin11),
    .sum(s51),
    .cout(c51)
);
Full_adder a61(
    .A(s51),
    .B(cin12),
    .cin(cin13),
    .sum(s61),
    .cout(c61)
);

endmodule

module adder4(
    input c0,
    input p0,
    input p1,
    input p2,
    input p3,
    input g0,
    input g1,
    input g2,
    input g3,
    output c1,
    output c2,
    output c3,
    output P,
    output G
);
assign c1 = g0 | p0&c0;
assign c2 = g1 | p1&g0 | p1&p0&c0;
assign c3 = g2 | p2&g1 | p2&p1&g0 | p2&p1&p0&c0;
assign P = p3&p2&p1&p0;
assign G = g3 | p3&g2 | p3&p2&g1 | p3&p2&p1&g0;

endmodule

module adder64(
    input cin,
    input [63:0] A,
    input [63:0] B,
    output [63:0] sum,
    output cout
);
wire p0_0,p0_1,p0_2,p0_3,p0_4,p0_5,p0_6,p0_7,p0_8,p0_9,p0_10,p0_11,p0_12,p0_13,p0_14,p0_15,p0_16,p0_17,p0_18,p0_19,p0_20,p0_21,p0_22,p0_23,p0_24,p0_25,p0_26,p0_27,p0_28,p0_29,p0_30,p0_31,p0_32,p0_33,p0_34,p0_35,p0_36,p0_37,p0_38,p0_39,p0_40,p0_41,p0_42,p0_43,p0_44,p0_45,p0_46,p0_47,p0_48,p0_49,p0_50,p0_51,p0_52,p0_53,p0_54,p0_55,p0_56,p0_57,p0_58,p0_59,p0_60,p0_61,p0_62,p0_63;
wire g0_0,g0_1,g0_2,g0_3,g0_4,g0_5,g0_6,g0_7,g0_8,g0_9,g0_10,g0_11,g0_12,g0_13,g0_14,g0_15,g0_16,g0_17,g0_18,g0_19,g0_20,g0_21,g0_22,g0_23,g0_24,g0_25,g0_26,g0_27,g0_28,g0_29,g0_30,g0_31,g0_32,g0_33,g0_34,g0_35,g0_36,g0_37,g0_38,g0_39,g0_40,g0_41,g0_42,g0_43,g0_44,g0_45,g0_46,g0_47,g0_48,g0_49,g0_50,g0_51,g0_52,g0_53,g0_54,g0_55,g0_56,g0_57,g0_58,g0_59,g0_60,g0_61,g0_62,g0_63;
wire c1_1,c1_2,c1_3,c1_5,c1_6,c1_7,c1_9,c1_10,c1_11,c1_13,c1_14,c1_15,c1_17,c1_18,c1_19,c1_21,c1_22,c1_23,c1_25,c1_26,c1_27,c1_29,c1_30,c1_31,c1_33,c1_34,c1_35,c1_37,c1_38,c1_39,c1_41,c1_42,c1_43,c1_45,c1_46,c1_47,c1_49,c1_50,c1_51,c1_53,c1_54,c1_55,c1_57,c1_58,c1_59,c1_61,c1_62,c1_63;
wire p1_0,p1_1,p1_2,p1_3,p1_5,p1_6,p1_7,p1_9,p1_10,p1_11,p1_13,p1_14,p1_15;
wire g1_0,g1_1,g1_2,g1_3,g1_5,g1_6,g1_7,g1_9,g1_10,g1_11,g1_13,g1_14,g1_15;
wire c2_1,c2_2,c2_3,c2_5,c2_6,c2_7,c2_9,c2_10,c2_11,c2_13,c2_14,c2_15;
wire p2_0,p2_1,p2_2,p2_3;
wire g2_0,g2_1,g2_2,g2_3;
wire c3_1,c3_2,c3_3;
wire p3_0,g3_0;

assign cout = p3_0 & cin | g3_0;

assign p0_0 = A[0] | B[0];
assign p0_1 = A[1] | B[1];
assign p0_2 = A[2] | B[2];
assign p0_3 = A[3] | B[3];
assign p0_4 = A[4] | B[4];
assign p0_5 = A[5] | B[5];
assign p0_6 = A[6] | B[6];
assign p0_7 = A[7] | B[7];
assign p0_8 = A[8] | B[8];
assign p0_9 = A[9] | B[9];
assign p0_10 = A[10] | B[10];
assign p0_11 = A[11] | B[11];
assign p0_12 = A[12] | B[12];
assign p0_13 = A[13] | B[13];
assign p0_14 = A[14] | B[14];
assign p0_15 = A[15] | B[15];
assign p0_16 = A[16] | B[16];
assign p0_17 = A[17] | B[17];
assign p0_18 = A[18] | B[18];
assign p0_19 = A[19] | B[19];
assign p0_20 = A[20] | B[20];
assign p0_21 = A[21] | B[21];
assign p0_22 = A[22] | B[22];
assign p0_23 = A[23] | B[23];
assign p0_24 = A[24] | B[24];
assign p0_25 = A[25] | B[25];
assign p0_26 = A[26] | B[26];
assign p0_27 = A[27] | B[27];
assign p0_28 = A[28] | B[28];
assign p0_29 = A[29] | B[29];
assign p0_30 = A[30] | B[30];
assign p0_31 = A[31] | B[31];
assign p0_32 = A[32] | B[32];
assign p0_33 = A[33] | B[33];
assign p0_34 = A[34] | B[34];
assign p0_35 = A[35] | B[35];
assign p0_36 = A[36] | B[36];
assign p0_37 = A[37] | B[37];
assign p0_38 = A[38] | B[38];
assign p0_39 = A[39] | B[39];
assign p0_40 = A[40] | B[40];
assign p0_41 = A[41] | B[41];
assign p0_42 = A[42] | B[42];
assign p0_43 = A[43] | B[43];
assign p0_44 = A[44] | B[44];
assign p0_45 = A[45] | B[45];
assign p0_46 = A[46] | B[46];
assign p0_47 = A[47] | B[47];
assign p0_48 = A[48] | B[48];
assign p0_49 = A[49] | B[49];
assign p0_50 = A[50] | B[50];
assign p0_51 = A[51] | B[51];
assign p0_52 = A[52] | B[52];
assign p0_53 = A[53] | B[53];
assign p0_54 = A[54] | B[54];
assign p0_55 = A[55] | B[55];
assign p0_56 = A[56] | B[56];
assign p0_57 = A[57] | B[57];
assign p0_58 = A[58] | B[58];
assign p0_59 = A[59] | B[59];
assign p0_60 = A[60] | B[60];
assign p0_61 = A[61] | B[61];
assign p0_62 = A[62] | B[62];
assign p0_63 = A[63] | B[63];
assign g0_0 = A[0] & B[0];
assign g0_1 = A[1] & B[1];
assign g0_2 = A[2] & B[2];
assign g0_3 = A[3] & B[3];
assign g0_4 = A[4] & B[4];
assign g0_5 = A[5] & B[5];
assign g0_6 = A[6] & B[6];
assign g0_7 = A[7] & B[7];
assign g0_8 = A[8] & B[8];
assign g0_9 = A[9] & B[9];
assign g0_10 = A[10] & B[10];
assign g0_11 = A[11] & B[11];
assign g0_12 = A[12] & B[12];
assign g0_13 = A[13] & B[13];
assign g0_14 = A[14] & B[14];
assign g0_15 = A[15] & B[15];
assign g0_16 = A[16] & B[16];
assign g0_17 = A[17] & B[17];
assign g0_18 = A[18] & B[18];
assign g0_19 = A[19] & B[19];
assign g0_20 = A[20] & B[20];
assign g0_21 = A[21] & B[21];
assign g0_22 = A[22] & B[22];
assign g0_23 = A[23] & B[23];
assign g0_24 = A[24] & B[24];
assign g0_25 = A[25] & B[25];
assign g0_26 = A[26] & B[26];
assign g0_27 = A[27] & B[27];
assign g0_28 = A[28] & B[28];
assign g0_29 = A[29] & B[29];
assign g0_30 = A[30] & B[30];
assign g0_31 = A[31] & B[31];
assign g0_32 = A[32] & B[32];
assign g0_33 = A[33] & B[33];
assign g0_34 = A[34] & B[34];
assign g0_35 = A[35] & B[35];
assign g0_36 = A[36] & B[36];
assign g0_37 = A[37] & B[37];
assign g0_38 = A[38] & B[38];
assign g0_39 = A[39] & B[39];
assign g0_40 = A[40] & B[40];
assign g0_41 = A[41] & B[41];
assign g0_42 = A[42] & B[42];
assign g0_43 = A[43] & B[43];
assign g0_44 = A[44] & B[44];
assign g0_45 = A[45] & B[45];
assign g0_46 = A[46] & B[46];
assign g0_47 = A[47] & B[47];
assign g0_48 = A[48] & B[48];
assign g0_49 = A[49] & B[49];
assign g0_50 = A[50] & B[50];
assign g0_51 = A[51] & B[51];
assign g0_52 = A[52] & B[52];
assign g0_53 = A[53] & B[53];
assign g0_54 = A[54] & B[54];
assign g0_55 = A[55] & B[55];
assign g0_56 = A[56] & B[56];
assign g0_57 = A[57] & B[57];
assign g0_58 = A[58] & B[58];
assign g0_59 = A[59] & B[59];
assign g0_60 = A[60] & B[60];
assign g0_61 = A[61] & B[61];
assign g0_62 = A[62] & B[62];
assign g0_63 = A[63] & B[63];

adder4 add1_0(
	.c0(cin),
	.p0(p0_0),
	.p1(p0_1),
	.p2(p0_2),
	.p3(p0_3),
	.g0(g0_0),
	.g1(g0_1),
	.g2(g0_2),
	.g3(g0_3),
	.c1(c1_1),
	.c2(c1_2),
	.c3(c1_3),
	.P(p1_0),
	.G(g1_0)
);
adder4 add1_1(
	.c0(c2_1),
	.p0(p0_4),
	.p1(p0_5),
	.p2(p0_6),
	.p3(p0_7),
	.g0(g0_4),
	.g1(g0_5),
	.g2(g0_6),
	.g3(g0_7),
	.c1(c1_5),
	.c2(c1_6),
	.c3(c1_7),
	.P(p1_1),
	.G(g1_1)
);
adder4 add1_2(
	.c0(c2_2),
	.p0(p0_8),
	.p1(p0_9),
	.p2(p0_10),
	.p3(p0_11),
	.g0(g0_8),
	.g1(g0_9),
	.g2(g0_10),
	.g3(g0_11),
	.c1(c1_9),
	.c2(c1_10),
	.c3(c1_11),
	.P(p1_2),
	.G(g1_2)
);
adder4 add1_3(
	.c0(c2_3),
	.p0(p0_12),
	.p1(p0_13),
	.p2(p0_14),
	.p3(p0_15),
	.g0(g0_12),
	.g1(g0_13),
	.g2(g0_14),
	.g3(g0_15),
	.c1(c1_13),
	.c2(c1_14),
	.c3(c1_15),
	.P(p1_3),
	.G(g1_3)
);
adder4 add1_4(
	.c0(c3_1),
	.p0(p0_16),
	.p1(p0_17),
	.p2(p0_18),
	.p3(p0_19),
	.g0(g0_16),
	.g1(g0_17),
	.g2(g0_18),
	.g3(g0_19),
	.c1(c1_17),
	.c2(c1_18),
	.c3(c1_19),
	.P(p1_4),
	.G(g1_4)
);
adder4 add1_5(
	.c0(c2_5),
	.p0(p0_20),
	.p1(p0_21),
	.p2(p0_22),
	.p3(p0_23),
	.g0(g0_20),
	.g1(g0_21),
	.g2(g0_22),
	.g3(g0_23),
	.c1(c1_21),
	.c2(c1_22),
	.c3(c1_23),
	.P(p1_5),
	.G(g1_5)
);
adder4 add1_6(
	.c0(c2_6),
	.p0(p0_24),
	.p1(p0_25),
	.p2(p0_26),
	.p3(p0_27),
	.g0(g0_24),
	.g1(g0_25),
	.g2(g0_26),
	.g3(g0_27),
	.c1(c1_25),
	.c2(c1_26),
	.c3(c1_27),
	.P(p1_6),
	.G(g1_6)
);
adder4 add1_7(
	.c0(c2_7),
	.p0(p0_28),
	.p1(p0_29),
	.p2(p0_30),
	.p3(p0_31),
	.g0(g0_28),
	.g1(g0_29),
	.g2(g0_30),
	.g3(g0_31),
	.c1(c1_29),
	.c2(c1_30),
	.c3(c1_31),
	.P(p1_7),
	.G(g1_7)
);
adder4 add1_8(
	.c0(c3_2),
	.p0(p0_32),
	.p1(p0_33),
	.p2(p0_34),
	.p3(p0_35),
	.g0(g0_32),
	.g1(g0_33),
	.g2(g0_34),
	.g3(g0_35),
	.c1(c1_33),
	.c2(c1_34),
	.c3(c1_35),
	.P(p1_8),
	.G(g1_8)
);
adder4 add1_9(
	.c0(c2_9),
	.p0(p0_36),
	.p1(p0_37),
	.p2(p0_38),
	.p3(p0_39),
	.g0(g0_36),
	.g1(g0_37),
	.g2(g0_38),
	.g3(g0_39),
	.c1(c1_37),
	.c2(c1_38),
	.c3(c1_39),
	.P(p1_9),
	.G(g1_9)
);
adder4 add1_10(
	.c0(c2_10),
	.p0(p0_40),
	.p1(p0_41),
	.p2(p0_42),
	.p3(p0_43),
	.g0(g0_40),
	.g1(g0_41),
	.g2(g0_42),
	.g3(g0_43),
	.c1(c1_41),
	.c2(c1_42),
	.c3(c1_43),
	.P(p1_10),
	.G(g1_10)
);
adder4 add1_11(
	.c0(c2_11),
	.p0(p0_44),
	.p1(p0_45),
	.p2(p0_46),
	.p3(p0_47),
	.g0(g0_44),
	.g1(g0_45),
	.g2(g0_46),
	.g3(g0_47),
	.c1(c1_45),
	.c2(c1_46),
	.c3(c1_47),
	.P(p1_11),
	.G(g1_11)
);
adder4 add1_12(
	.c0(c3_3),
	.p0(p0_48),
	.p1(p0_49),
	.p2(p0_50),
	.p3(p0_51),
	.g0(g0_48),
	.g1(g0_49),
	.g2(g0_50),
	.g3(g0_51),
	.c1(c1_49),
	.c2(c1_50),
	.c3(c1_51),
	.P(p1_12),
	.G(g1_12)
);
adder4 add1_13(
	.c0(c2_13),
	.p0(p0_52),
	.p1(p0_53),
	.p2(p0_54),
	.p3(p0_55),
	.g0(g0_52),
	.g1(g0_53),
	.g2(g0_54),
	.g3(g0_55),
	.c1(c1_53),
	.c2(c1_54),
	.c3(c1_55),
	.P(p1_13),
	.G(g1_13)
);
adder4 add1_14(
	.c0(c2_14),
	.p0(p0_56),
	.p1(p0_57),
	.p2(p0_58),
	.p3(p0_59),
	.g0(g0_56),
	.g1(g0_57),
	.g2(g0_58),
	.g3(g0_59),
	.c1(c1_57),
	.c2(c1_58),
	.c3(c1_59),
	.P(p1_14),
	.G(g1_14)
);
adder4 add1_15(
	.c0(c2_15),
	.p0(p0_60),
	.p1(p0_61),
	.p2(p0_62),
	.p3(p0_63),
	.g0(g0_60),
	.g1(g0_61),
	.g2(g0_62),
	.g3(g0_63),
	.c1(c1_61),
	.c2(c1_62),
	.c3(c1_63),
	.P(p1_15),
	.G(g1_15)
);
adder4 add2_0(
	.c0(cin),
	.p0(p1_0),
	.p1(p1_1),
	.p2(p1_2),
	.p3(p1_3),
	.g0(g1_0),
	.g1(g1_1),
	.g2(g1_2),
	.g3(g1_3),
	.c1(c2_1),
	.c2(c2_2),
	.c3(c2_3),
	.P(p2_0),
	.G(g2_0)
);
adder4 add2_1(
	.c0(c3_1),
	.p0(p1_4),
	.p1(p1_5),
	.p2(p1_6),
	.p3(p1_7),
	.g0(g1_4),
	.g1(g1_5),
	.g2(g1_6),
	.g3(g1_7),
	.c1(c2_5),
	.c2(c2_6),
	.c3(c2_7),
	.P(p2_1),
	.G(g2_1)
);
adder4 add2_2(
	.c0(c3_2),
	.p0(p1_8),
	.p1(p1_9),
	.p2(p1_10),
	.p3(p1_11),
	.g0(g1_8),
	.g1(g1_9),
	.g2(g1_10),
	.g3(g1_11),
	.c1(c2_9),
	.c2(c2_10),
	.c3(c2_11),
	.P(p2_2),
	.G(g2_2)
);
adder4 add2_3(
	.c0(c3_3),
	.p0(p1_12),
	.p1(p1_13),
	.p2(p1_14),
	.p3(p1_15),
	.g0(g1_12),
	.g1(g1_13),
	.g2(g1_14),
	.g3(g1_15),
	.c1(c2_13),
	.c2(c2_14),
	.c3(c2_15),
	.P(p2_3),
	.G(g2_3)
);
adder4 add3_0(
	.c0(cin),
	.p0(p2_0),
	.p1(p2_1),
	.p2(p2_2),
	.p3(p2_3),
	.g0(g2_0),
	.g1(g2_1),
	.g2(g2_2),
	.g3(g2_3),
	.c1(c3_1),
	.c2(c3_2),
	.c3(c3_3),
	.P(p3_0),
	.G(g3_0)
);
Full_adder fa0(
	.A(A[0]),
	.B(B[0]),
	.cin(cin),
	.sum(sum[0]),
	.cout()
);
Full_adder fa1(
	.A(A[1]),
	.B(B[1]),
	.cin(c1_1),
	.sum(sum[1]),
	.cout()
);
Full_adder fa2(
	.A(A[2]),
	.B(B[2]),
	.cin(c1_2),
	.sum(sum[2]),
	.cout()
);
Full_adder fa3(
	.A(A[3]),
	.B(B[3]),
	.cin(c1_3),
	.sum(sum[3]),
	.cout()
);
Full_adder fa4(
	.A(A[4]),
	.B(B[4]),
	.cin(c2_1),
	.sum(sum[4]),
	.cout()
);
Full_adder fa5(
	.A(A[5]),
	.B(B[5]),
	.cin(c1_5),
	.sum(sum[5]),
	.cout()
);
Full_adder fa6(
	.A(A[6]),
	.B(B[6]),
	.cin(c1_6),
	.sum(sum[6]),
	.cout()
);
Full_adder fa7(
	.A(A[7]),
	.B(B[7]),
	.cin(c1_7),
	.sum(sum[7]),
	.cout()
);
Full_adder fa8(
	.A(A[8]),
	.B(B[8]),
	.cin(c2_2),
	.sum(sum[8]),
	.cout()
);
Full_adder fa9(
	.A(A[9]),
	.B(B[9]),
	.cin(c1_9),
	.sum(sum[9]),
	.cout()
);
Full_adder fa10(
	.A(A[10]),
	.B(B[10]),
	.cin(c1_10),
	.sum(sum[10]),
	.cout()
);
Full_adder fa11(
	.A(A[11]),
	.B(B[11]),
	.cin(c1_11),
	.sum(sum[11]),
	.cout()
);
Full_adder fa12(
	.A(A[12]),
	.B(B[12]),
	.cin(c2_3),
	.sum(sum[12]),
	.cout()
);
Full_adder fa13(
	.A(A[13]),
	.B(B[13]),
	.cin(c1_13),
	.sum(sum[13]),
	.cout()
);
Full_adder fa14(
	.A(A[14]),
	.B(B[14]),
	.cin(c1_14),
	.sum(sum[14]),
	.cout()
);
Full_adder fa15(
	.A(A[15]),
	.B(B[15]),
	.cin(c1_15),
	.sum(sum[15]),
	.cout()
);
Full_adder fa16(
	.A(A[16]),
	.B(B[16]),
	.cin(c3_1),
	.sum(sum[16]),
	.cout()
);
Full_adder fa17(
	.A(A[17]),
	.B(B[17]),
	.cin(c1_17),
	.sum(sum[17]),
	.cout()
);
Full_adder fa18(
	.A(A[18]),
	.B(B[18]),
	.cin(c1_18),
	.sum(sum[18]),
	.cout()
);
Full_adder fa19(
	.A(A[19]),
	.B(B[19]),
	.cin(c1_19),
	.sum(sum[19]),
	.cout()
);
Full_adder fa20(
	.A(A[20]),
	.B(B[20]),
	.cin(c2_5),
	.sum(sum[20]),
	.cout()
);
Full_adder fa21(
	.A(A[21]),
	.B(B[21]),
	.cin(c1_21),
	.sum(sum[21]),
	.cout()
);
Full_adder fa22(
	.A(A[22]),
	.B(B[22]),
	.cin(c1_22),
	.sum(sum[22]),
	.cout()
);
Full_adder fa23(
	.A(A[23]),
	.B(B[23]),
	.cin(c1_23),
	.sum(sum[23]),
	.cout()
);
Full_adder fa24(
	.A(A[24]),
	.B(B[24]),
	.cin(c2_6),
	.sum(sum[24]),
	.cout()
);
Full_adder fa25(
	.A(A[25]),
	.B(B[25]),
	.cin(c1_25),
	.sum(sum[25]),
	.cout()
);
Full_adder fa26(
	.A(A[26]),
	.B(B[26]),
	.cin(c1_26),
	.sum(sum[26]),
	.cout()
);
Full_adder fa27(
	.A(A[27]),
	.B(B[27]),
	.cin(c1_27),
	.sum(sum[27]),
	.cout()
);
Full_adder fa28(
	.A(A[28]),
	.B(B[28]),
	.cin(c2_7),
	.sum(sum[28]),
	.cout()
);
Full_adder fa29(
	.A(A[29]),
	.B(B[29]),
	.cin(c1_29),
	.sum(sum[29]),
	.cout()
);
Full_adder fa30(
	.A(A[30]),
	.B(B[30]),
	.cin(c1_30),
	.sum(sum[30]),
	.cout()
);
Full_adder fa31(
	.A(A[31]),
	.B(B[31]),
	.cin(c1_31),
	.sum(sum[31]),
	.cout()
);
Full_adder fa32(
	.A(A[32]),
	.B(B[32]),
	.cin(c3_2),
	.sum(sum[32]),
	.cout()
);
Full_adder fa33(
	.A(A[33]),
	.B(B[33]),
	.cin(c1_33),
	.sum(sum[33]),
	.cout()
);
Full_adder fa34(
	.A(A[34]),
	.B(B[34]),
	.cin(c1_34),
	.sum(sum[34]),
	.cout()
);
Full_adder fa35(
	.A(A[35]),
	.B(B[35]),
	.cin(c1_35),
	.sum(sum[35]),
	.cout()
);
Full_adder fa36(
	.A(A[36]),
	.B(B[36]),
	.cin(c2_9),
	.sum(sum[36]),
	.cout()
);
Full_adder fa37(
	.A(A[37]),
	.B(B[37]),
	.cin(c1_37),
	.sum(sum[37]),
	.cout()
);
Full_adder fa38(
	.A(A[38]),
	.B(B[38]),
	.cin(c1_38),
	.sum(sum[38]),
	.cout()
);
Full_adder fa39(
	.A(A[39]),
	.B(B[39]),
	.cin(c1_39),
	.sum(sum[39]),
	.cout()
);
Full_adder fa40(
	.A(A[40]),
	.B(B[40]),
	.cin(c2_10),
	.sum(sum[40]),
	.cout()
);
Full_adder fa41(
	.A(A[41]),
	.B(B[41]),
	.cin(c1_41),
	.sum(sum[41]),
	.cout()
);
Full_adder fa42(
	.A(A[42]),
	.B(B[42]),
	.cin(c1_42),
	.sum(sum[42]),
	.cout()
);
Full_adder fa43(
	.A(A[43]),
	.B(B[43]),
	.cin(c1_43),
	.sum(sum[43]),
	.cout()
);
Full_adder fa44(
	.A(A[44]),
	.B(B[44]),
	.cin(c2_11),
	.sum(sum[44]),
	.cout()
);
Full_adder fa45(
	.A(A[45]),
	.B(B[45]),
	.cin(c1_45),
	.sum(sum[45]),
	.cout()
);
Full_adder fa46(
	.A(A[46]),
	.B(B[46]),
	.cin(c1_46),
	.sum(sum[46]),
	.cout()
);
Full_adder fa47(
	.A(A[47]),
	.B(B[47]),
	.cin(c1_47),
	.sum(sum[47]),
	.cout()
);
Full_adder fa48(
	.A(A[48]),
	.B(B[48]),
	.cin(c3_3),
	.sum(sum[48]),
	.cout()
);
Full_adder fa49(
	.A(A[49]),
	.B(B[49]),
	.cin(c1_49),
	.sum(sum[49]),
	.cout()
);
Full_adder fa50(
	.A(A[50]),
	.B(B[50]),
	.cin(c1_50),
	.sum(sum[50]),
	.cout()
);
Full_adder fa51(
	.A(A[51]),
	.B(B[51]),
	.cin(c1_51),
	.sum(sum[51]),
	.cout()
);
Full_adder fa52(
	.A(A[52]),
	.B(B[52]),
	.cin(c2_13),
	.sum(sum[52]),
	.cout()
);
Full_adder fa53(
	.A(A[53]),
	.B(B[53]),
	.cin(c1_53),
	.sum(sum[53]),
	.cout()
);
Full_adder fa54(
	.A(A[54]),
	.B(B[54]),
	.cin(c1_54),
	.sum(sum[54]),
	.cout()
);
Full_adder fa55(
	.A(A[55]),
	.B(B[55]),
	.cin(c1_55),
	.sum(sum[55]),
	.cout()
);
Full_adder fa56(
	.A(A[56]),
	.B(B[56]),
	.cin(c2_14),
	.sum(sum[56]),
	.cout()
);
Full_adder fa57(
	.A(A[57]),
	.B(B[57]),
	.cin(c1_57),
	.sum(sum[57]),
	.cout()
);
Full_adder fa58(
	.A(A[58]),
	.B(B[58]),
	.cin(c1_58),
	.sum(sum[58]),
	.cout()
);
Full_adder fa59(
	.A(A[59]),
	.B(B[59]),
	.cin(c1_59),
	.sum(sum[59]),
	.cout()
);
Full_adder fa60(
	.A(A[60]),
	.B(B[60]),
	.cin(c2_15),
	.sum(sum[60]),
	.cout()
);
Full_adder fa61(
	.A(A[61]),
	.B(B[61]),
	.cin(c1_61),
	.sum(sum[61]),
	.cout()
);
Full_adder fa62(
	.A(A[62]),
	.B(B[62]),
	.cin(c1_62),
	.sum(sum[62]),
	.cout()
);
Full_adder fa63(
	.A(A[63]),
	.B(B[63]),
	.cin(c1_63),
	.sum(sum[63]),
	.cout()
);


endmodule


